// This is the unpowered netlist.
module RAM32_1RW1R (CLK,
    EN0,
    EN1,
    A0,
    A1,
    Di0,
    Do0,
    Do1,
    WE0);
 input CLK;
 input EN0;
 input EN1;
 input [4:0] A0;
 input [4:0] A1;
 input [31:0] Di0;
 output [31:0] Do0;
 output [31:0] Do1;
 input [3:0] WE0;

 wire \A0BUF[0].X ;
 wire \A0BUF[1].X ;
 wire \A0BUF[2].X ;
 wire \A0BUF[3].X ;
 wire \A0BUF[4].X ;
 wire \A1BUF[0].X ;
 wire \A1BUF[1].X ;
 wire \A1BUF[2].X ;
 wire \A1BUF[3].X ;
 wire \A1BUF[4].X ;
 wire \BYTE[0].FLOATBUF0[0].A ;
 wire \BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BYTE[0].FLOATBUF0[0].TE_BN ;
 wire \BYTE[0].FLOATBUF0[0].Z ;
 wire \BYTE[0].FLOATBUF0[1].TE_BN ;
 wire \BYTE[0].FLOATBUF0[1].Z ;
 wire \BYTE[0].FLOATBUF0[2].TE_BN ;
 wire \BYTE[0].FLOATBUF0[2].Z ;
 wire \BYTE[0].FLOATBUF0[3].TE_BN ;
 wire \BYTE[0].FLOATBUF0[3].Z ;
 wire \BYTE[0].FLOATBUF0[4].TE_BN ;
 wire \BYTE[0].FLOATBUF0[4].Z ;
 wire \BYTE[0].FLOATBUF0[5].TE_BN ;
 wire \BYTE[0].FLOATBUF0[5].Z ;
 wire \BYTE[0].FLOATBUF0[6].TE_BN ;
 wire \BYTE[0].FLOATBUF0[6].Z ;
 wire \BYTE[0].FLOATBUF0[7].TE_BN ;
 wire \BYTE[0].FLOATBUF0[7].Z ;
 wire \BYTE[0].FLOATBUF1[0].A ;
 wire \BYTE[0].FLOATBUF1[0].TE_B ;
 wire \BYTE[0].FLOATBUF1[0].TE_BN ;
 wire \BYTE[0].FLOATBUF1[0].Z ;
 wire \BYTE[0].FLOATBUF1[1].TE_BN ;
 wire \BYTE[0].FLOATBUF1[1].Z ;
 wire \BYTE[0].FLOATBUF1[2].TE_BN ;
 wire \BYTE[0].FLOATBUF1[2].Z ;
 wire \BYTE[0].FLOATBUF1[3].TE_BN ;
 wire \BYTE[0].FLOATBUF1[3].Z ;
 wire \BYTE[0].FLOATBUF1[4].TE_BN ;
 wire \BYTE[0].FLOATBUF1[4].Z ;
 wire \BYTE[0].FLOATBUF1[5].TE_BN ;
 wire \BYTE[0].FLOATBUF1[5].Z ;
 wire \BYTE[0].FLOATBUF1[6].TE_BN ;
 wire \BYTE[0].FLOATBUF1[6].Z ;
 wire \BYTE[0].FLOATBUF1[7].TE_BN ;
 wire \BYTE[0].FLOATBUF1[7].Z ;
 wire \BYTE[1].FLOATBUF0[10].A ;
 wire \BYTE[1].FLOATBUF0[10].TE_B ;
 wire \BYTE[1].FLOATBUF0[10].TE_BN ;
 wire \BYTE[1].FLOATBUF0[10].Z ;
 wire \BYTE[1].FLOATBUF0[11].TE_BN ;
 wire \BYTE[1].FLOATBUF0[11].Z ;
 wire \BYTE[1].FLOATBUF0[12].TE_BN ;
 wire \BYTE[1].FLOATBUF0[12].Z ;
 wire \BYTE[1].FLOATBUF0[13].TE_BN ;
 wire \BYTE[1].FLOATBUF0[13].Z ;
 wire \BYTE[1].FLOATBUF0[14].TE_BN ;
 wire \BYTE[1].FLOATBUF0[14].Z ;
 wire \BYTE[1].FLOATBUF0[15].TE_BN ;
 wire \BYTE[1].FLOATBUF0[15].Z ;
 wire \BYTE[1].FLOATBUF0[8].TE_BN ;
 wire \BYTE[1].FLOATBUF0[8].Z ;
 wire \BYTE[1].FLOATBUF0[9].TE_BN ;
 wire \BYTE[1].FLOATBUF0[9].Z ;
 wire \BYTE[1].FLOATBUF1[10].A ;
 wire \BYTE[1].FLOATBUF1[10].TE_B ;
 wire \BYTE[1].FLOATBUF1[10].TE_BN ;
 wire \BYTE[1].FLOATBUF1[10].Z ;
 wire \BYTE[1].FLOATBUF1[11].TE_BN ;
 wire \BYTE[1].FLOATBUF1[11].Z ;
 wire \BYTE[1].FLOATBUF1[12].TE_BN ;
 wire \BYTE[1].FLOATBUF1[12].Z ;
 wire \BYTE[1].FLOATBUF1[13].TE_BN ;
 wire \BYTE[1].FLOATBUF1[13].Z ;
 wire \BYTE[1].FLOATBUF1[14].TE_BN ;
 wire \BYTE[1].FLOATBUF1[14].Z ;
 wire \BYTE[1].FLOATBUF1[15].TE_BN ;
 wire \BYTE[1].FLOATBUF1[15].Z ;
 wire \BYTE[1].FLOATBUF1[8].TE_BN ;
 wire \BYTE[1].FLOATBUF1[8].Z ;
 wire \BYTE[1].FLOATBUF1[9].TE_BN ;
 wire \BYTE[1].FLOATBUF1[9].Z ;
 wire \BYTE[2].FLOATBUF0[16].A ;
 wire \BYTE[2].FLOATBUF0[16].TE_B ;
 wire \BYTE[2].FLOATBUF0[16].TE_BN ;
 wire \BYTE[2].FLOATBUF0[16].Z ;
 wire \BYTE[2].FLOATBUF0[17].TE_BN ;
 wire \BYTE[2].FLOATBUF0[17].Z ;
 wire \BYTE[2].FLOATBUF0[18].TE_BN ;
 wire \BYTE[2].FLOATBUF0[18].Z ;
 wire \BYTE[2].FLOATBUF0[19].TE_BN ;
 wire \BYTE[2].FLOATBUF0[19].Z ;
 wire \BYTE[2].FLOATBUF0[20].TE_BN ;
 wire \BYTE[2].FLOATBUF0[20].Z ;
 wire \BYTE[2].FLOATBUF0[21].TE_BN ;
 wire \BYTE[2].FLOATBUF0[21].Z ;
 wire \BYTE[2].FLOATBUF0[22].TE_BN ;
 wire \BYTE[2].FLOATBUF0[22].Z ;
 wire \BYTE[2].FLOATBUF0[23].TE_BN ;
 wire \BYTE[2].FLOATBUF0[23].Z ;
 wire \BYTE[2].FLOATBUF1[16].A ;
 wire \BYTE[2].FLOATBUF1[16].TE_B ;
 wire \BYTE[2].FLOATBUF1[16].TE_BN ;
 wire \BYTE[2].FLOATBUF1[16].Z ;
 wire \BYTE[2].FLOATBUF1[17].TE_BN ;
 wire \BYTE[2].FLOATBUF1[17].Z ;
 wire \BYTE[2].FLOATBUF1[18].TE_BN ;
 wire \BYTE[2].FLOATBUF1[18].Z ;
 wire \BYTE[2].FLOATBUF1[19].TE_BN ;
 wire \BYTE[2].FLOATBUF1[19].Z ;
 wire \BYTE[2].FLOATBUF1[20].TE_BN ;
 wire \BYTE[2].FLOATBUF1[20].Z ;
 wire \BYTE[2].FLOATBUF1[21].TE_BN ;
 wire \BYTE[2].FLOATBUF1[21].Z ;
 wire \BYTE[2].FLOATBUF1[22].TE_BN ;
 wire \BYTE[2].FLOATBUF1[22].Z ;
 wire \BYTE[2].FLOATBUF1[23].TE_BN ;
 wire \BYTE[2].FLOATBUF1[23].Z ;
 wire \BYTE[3].FLOATBUF0[24].A ;
 wire \BYTE[3].FLOATBUF0[24].TE_B ;
 wire \BYTE[3].FLOATBUF0[24].TE_BN ;
 wire \BYTE[3].FLOATBUF0[24].Z ;
 wire \BYTE[3].FLOATBUF0[25].TE_BN ;
 wire \BYTE[3].FLOATBUF0[25].Z ;
 wire \BYTE[3].FLOATBUF0[26].TE_BN ;
 wire \BYTE[3].FLOATBUF0[26].Z ;
 wire \BYTE[3].FLOATBUF0[27].TE_BN ;
 wire \BYTE[3].FLOATBUF0[27].Z ;
 wire \BYTE[3].FLOATBUF0[28].TE_BN ;
 wire \BYTE[3].FLOATBUF0[28].Z ;
 wire \BYTE[3].FLOATBUF0[29].TE_BN ;
 wire \BYTE[3].FLOATBUF0[29].Z ;
 wire \BYTE[3].FLOATBUF0[30].TE_BN ;
 wire \BYTE[3].FLOATBUF0[30].Z ;
 wire \BYTE[3].FLOATBUF0[31].TE_BN ;
 wire \BYTE[3].FLOATBUF0[31].Z ;
 wire \BYTE[3].FLOATBUF1[24].A ;
 wire \BYTE[3].FLOATBUF1[24].TE_B ;
 wire \BYTE[3].FLOATBUF1[24].TE_BN ;
 wire \BYTE[3].FLOATBUF1[24].Z ;
 wire \BYTE[3].FLOATBUF1[25].TE_BN ;
 wire \BYTE[3].FLOATBUF1[25].Z ;
 wire \BYTE[3].FLOATBUF1[26].TE_BN ;
 wire \BYTE[3].FLOATBUF1[26].Z ;
 wire \BYTE[3].FLOATBUF1[27].TE_BN ;
 wire \BYTE[3].FLOATBUF1[27].Z ;
 wire \BYTE[3].FLOATBUF1[28].TE_BN ;
 wire \BYTE[3].FLOATBUF1[28].Z ;
 wire \BYTE[3].FLOATBUF1[29].TE_BN ;
 wire \BYTE[3].FLOATBUF1[29].Z ;
 wire \BYTE[3].FLOATBUF1[30].TE_BN ;
 wire \BYTE[3].FLOATBUF1[30].Z ;
 wire \BYTE[3].FLOATBUF1[31].TE_BN ;
 wire \BYTE[3].FLOATBUF1[31].Z ;
 wire \CLKBUF.X ;
 wire \DEC0.A_N[0] ;
 wire \DEC0.A_N[1] ;
 wire \DEC0.EN ;
 wire \DEC0.EN_N ;
 wire \DEC1.A_N[0] ;
 wire \DEC1.A_N[1] ;
 wire \DEC1.EN ;
 wire \DEC1.EN_N ;
 wire \DIBUF[0].X ;
 wire \DIBUF[10].X ;
 wire \DIBUF[11].X ;
 wire \DIBUF[12].X ;
 wire \DIBUF[13].X ;
 wire \DIBUF[14].X ;
 wire \DIBUF[15].X ;
 wire \DIBUF[16].X ;
 wire \DIBUF[17].X ;
 wire \DIBUF[18].X ;
 wire \DIBUF[19].X ;
 wire \DIBUF[1].X ;
 wire \DIBUF[20].X ;
 wire \DIBUF[21].X ;
 wire \DIBUF[22].X ;
 wire \DIBUF[23].X ;
 wire \DIBUF[24].X ;
 wire \DIBUF[25].X ;
 wire \DIBUF[26].X ;
 wire \DIBUF[27].X ;
 wire \DIBUF[28].X ;
 wire \DIBUF[29].X ;
 wire \DIBUF[2].X ;
 wire \DIBUF[30].X ;
 wire \DIBUF[31].X ;
 wire \DIBUF[3].X ;
 wire \DIBUF[4].X ;
 wire \DIBUF[5].X ;
 wire \DIBUF[6].X ;
 wire \DIBUF[7].X ;
 wire \DIBUF[8].X ;
 wire \DIBUF[9].X ;
 wire \Do0_REG.CLKBUF[0] ;
 wire \Do0_REG.CLKBUF[1] ;
 wire \Do0_REG.CLKBUF[2] ;
 wire \Do0_REG.CLKBUF[3] ;
 wire \Do0_REG.CLK_buf ;
 wire \Do1_REG.CLKBUF[0] ;
 wire \Do1_REG.CLKBUF[1] ;
 wire \Do1_REG.CLKBUF[2] ;
 wire \Do1_REG.CLKBUF[3] ;
 wire \Do1_REG.CLK_buf ;
 wire \SLICE[0].RAM8.CLKBUF.X ;
 wire \SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[0].RAM8.DEC0.A_buf_N[0] ;
 wire \SLICE[0].RAM8.DEC0.A_buf_N[1] ;
 wire \SLICE[0].RAM8.DEC0.EN ;
 wire \SLICE[0].RAM8.DEC0.EN_buf ;
 wire \SLICE[0].RAM8.DEC0.EN_buf_N ;
 wire \SLICE[0].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[0].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[0].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[0].RAM8.DEC1.A_buf_N[0] ;
 wire \SLICE[0].RAM8.DEC1.A_buf_N[1] ;
 wire \SLICE[0].RAM8.DEC1.EN ;
 wire \SLICE[0].RAM8.DEC1.EN_buf ;
 wire \SLICE[0].RAM8.DEC1.EN_buf_N ;
 wire \SLICE[0].RAM8.WEBUF[0].A ;
 wire \SLICE[0].RAM8.WEBUF[0].X ;
 wire \SLICE[0].RAM8.WEBUF[1].A ;
 wire \SLICE[0].RAM8.WEBUF[1].X ;
 wire \SLICE[0].RAM8.WEBUF[2].A ;
 wire \SLICE[0].RAM8.WEBUF[2].X ;
 wire \SLICE[0].RAM8.WEBUF[3].A ;
 wire \SLICE[0].RAM8.WEBUF[3].X ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[1].RAM8.CLKBUF.X ;
 wire \SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[1].RAM8.DEC0.A_buf_N[0] ;
 wire \SLICE[1].RAM8.DEC0.A_buf_N[1] ;
 wire \SLICE[1].RAM8.DEC0.EN ;
 wire \SLICE[1].RAM8.DEC0.EN_buf ;
 wire \SLICE[1].RAM8.DEC0.EN_buf_N ;
 wire \SLICE[1].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[1].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[1].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[1].RAM8.DEC1.A_buf_N[0] ;
 wire \SLICE[1].RAM8.DEC1.A_buf_N[1] ;
 wire \SLICE[1].RAM8.DEC1.EN ;
 wire \SLICE[1].RAM8.DEC1.EN_buf ;
 wire \SLICE[1].RAM8.DEC1.EN_buf_N ;
 wire \SLICE[1].RAM8.WEBUF[0].X ;
 wire \SLICE[1].RAM8.WEBUF[1].X ;
 wire \SLICE[1].RAM8.WEBUF[2].X ;
 wire \SLICE[1].RAM8.WEBUF[3].X ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[2].RAM8.CLKBUF.X ;
 wire \SLICE[2].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[2].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[2].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[2].RAM8.DEC0.A_buf_N[0] ;
 wire \SLICE[2].RAM8.DEC0.A_buf_N[1] ;
 wire \SLICE[2].RAM8.DEC0.EN ;
 wire \SLICE[2].RAM8.DEC0.EN_buf ;
 wire \SLICE[2].RAM8.DEC0.EN_buf_N ;
 wire \SLICE[2].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[2].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[2].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[2].RAM8.DEC1.A_buf_N[0] ;
 wire \SLICE[2].RAM8.DEC1.A_buf_N[1] ;
 wire \SLICE[2].RAM8.DEC1.EN ;
 wire \SLICE[2].RAM8.DEC1.EN_buf ;
 wire \SLICE[2].RAM8.DEC1.EN_buf_N ;
 wire \SLICE[2].RAM8.WEBUF[0].X ;
 wire \SLICE[2].RAM8.WEBUF[1].X ;
 wire \SLICE[2].RAM8.WEBUF[2].X ;
 wire \SLICE[2].RAM8.WEBUF[3].X ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[3].RAM8.CLKBUF.X ;
 wire \SLICE[3].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[3].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[3].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[3].RAM8.DEC0.A_buf_N[0] ;
 wire \SLICE[3].RAM8.DEC0.A_buf_N[1] ;
 wire \SLICE[3].RAM8.DEC0.EN ;
 wire \SLICE[3].RAM8.DEC0.EN_buf ;
 wire \SLICE[3].RAM8.DEC0.EN_buf_N ;
 wire \SLICE[3].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[3].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[3].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[3].RAM8.DEC1.A_buf_N[0] ;
 wire \SLICE[3].RAM8.DEC1.A_buf_N[1] ;
 wire \SLICE[3].RAM8.DEC1.EN ;
 wire \SLICE[3].RAM8.DEC1.EN_buf ;
 wire \SLICE[3].RAM8.DEC1.EN_buf_N ;
 wire \SLICE[3].RAM8.WEBUF[0].X ;
 wire \SLICE[3].RAM8.WEBUF[1].X ;
 wire \SLICE[3].RAM8.WEBUF[2].X ;
 wire \SLICE[3].RAM8.WEBUF[3].X ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[7].W.SEL1 ;
 wire zero_;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[0].__cell__  (.I(A0[0]),
    .Z(\A0BUF[0].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[1].__cell__  (.I(A0[1]),
    .Z(\A0BUF[1].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[2].__cell__  (.I(A0[2]),
    .Z(\A0BUF[2].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[3].__cell__  (.I(A0[3]),
    .Z(\A0BUF[3].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[4].__cell__  (.I(A0[4]),
    .Z(\A0BUF[4].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[0].__cell__  (.I(A1[0]),
    .Z(\A1BUF[0].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[1].__cell__  (.I(A1[1]),
    .Z(\A1BUF[1].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[2].__cell__  (.I(A1[2]),
    .Z(\A1BUF[2].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[3].__cell__  (.I(A1[3]),
    .Z(\A1BUF[3].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[4].__cell__  (.I(A1[4]),
    .Z(\A1BUF[4].X ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[0].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[0].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[0].__cell__  (.EN(\BYTE[0].FLOATBUF0[0].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[1].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[1].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[1].__cell__  (.EN(\BYTE[0].FLOATBUF0[1].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[2].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[2].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[2].__cell__  (.EN(\BYTE[0].FLOATBUF0[2].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[3].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[3].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[3].__cell__  (.EN(\BYTE[0].FLOATBUF0[3].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[4].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[4].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[4].__cell__  (.EN(\BYTE[0].FLOATBUF0[4].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[5].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[5].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[5].__cell__  (.EN(\BYTE[0].FLOATBUF0[5].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[6].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[6].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[6].__cell__  (.EN(\BYTE[0].FLOATBUF0[6].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[7].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[7].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[7].__cell__  (.EN(\BYTE[0].FLOATBUF0[7].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[0].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[0].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[0].__cell__  (.EN(\BYTE[0].FLOATBUF1[0].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[1].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[1].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[1].__cell__  (.EN(\BYTE[0].FLOATBUF1[1].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[2].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[2].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[2].__cell__  (.EN(\BYTE[0].FLOATBUF1[2].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[3].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[3].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[3].__cell__  (.EN(\BYTE[0].FLOATBUF1[3].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[4].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[4].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[4].__cell__  (.EN(\BYTE[0].FLOATBUF1[4].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[5].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[5].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[5].__cell__  (.EN(\BYTE[0].FLOATBUF1[5].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[6].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[6].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[6].__cell__  (.EN(\BYTE[0].FLOATBUF1[6].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[7].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[7].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[7].__cell__  (.EN(\BYTE[0].FLOATBUF1[7].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[10].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[10].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[10].__cell__  (.EN(\BYTE[1].FLOATBUF0[10].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[11].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[11].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[11].__cell__  (.EN(\BYTE[1].FLOATBUF0[11].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[12].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[12].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[12].__cell__  (.EN(\BYTE[1].FLOATBUF0[12].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[13].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[13].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[13].__cell__  (.EN(\BYTE[1].FLOATBUF0[13].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[14].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[14].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[14].__cell__  (.EN(\BYTE[1].FLOATBUF0[14].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[15].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[15].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[15].__cell__  (.EN(\BYTE[1].FLOATBUF0[15].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[8].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[8].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[8].__cell__  (.EN(\BYTE[1].FLOATBUF0[8].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[9].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[9].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[9].__cell__  (.EN(\BYTE[1].FLOATBUF0[9].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[10].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[10].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[10].__cell__  (.EN(\BYTE[1].FLOATBUF1[10].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[11].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[11].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[11].__cell__  (.EN(\BYTE[1].FLOATBUF1[11].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[12].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[12].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[12].__cell__  (.EN(\BYTE[1].FLOATBUF1[12].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[13].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[13].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[13].__cell__  (.EN(\BYTE[1].FLOATBUF1[13].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[14].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[14].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[14].__cell__  (.EN(\BYTE[1].FLOATBUF1[14].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[15].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[15].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[15].__cell__  (.EN(\BYTE[1].FLOATBUF1[15].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[8].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[8].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[8].__cell__  (.EN(\BYTE[1].FLOATBUF1[8].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[9].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[9].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[9].__cell__  (.EN(\BYTE[1].FLOATBUF1[9].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[16].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[16].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[16].__cell__  (.EN(\BYTE[2].FLOATBUF0[16].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[17].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[17].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[17].__cell__  (.EN(\BYTE[2].FLOATBUF0[17].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[18].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[18].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[18].__cell__  (.EN(\BYTE[2].FLOATBUF0[18].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[19].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[19].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[19].__cell__  (.EN(\BYTE[2].FLOATBUF0[19].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[20].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[20].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[20].__cell__  (.EN(\BYTE[2].FLOATBUF0[20].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[21].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[21].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[21].__cell__  (.EN(\BYTE[2].FLOATBUF0[21].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[22].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[22].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[22].__cell__  (.EN(\BYTE[2].FLOATBUF0[22].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[23].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[23].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[23].__cell__  (.EN(\BYTE[2].FLOATBUF0[23].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[16].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[16].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[16].__cell__  (.EN(\BYTE[2].FLOATBUF1[16].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[17].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[17].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[17].__cell__  (.EN(\BYTE[2].FLOATBUF1[17].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[18].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[18].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[18].__cell__  (.EN(\BYTE[2].FLOATBUF1[18].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[19].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[19].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[19].__cell__  (.EN(\BYTE[2].FLOATBUF1[19].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[20].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[20].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[20].__cell__  (.EN(\BYTE[2].FLOATBUF1[20].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[21].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[21].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[21].__cell__  (.EN(\BYTE[2].FLOATBUF1[21].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[22].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[22].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[22].__cell__  (.EN(\BYTE[2].FLOATBUF1[22].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[23].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[23].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[23].__cell__  (.EN(\BYTE[2].FLOATBUF1[23].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[24].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[24].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[24].__cell__  (.EN(\BYTE[3].FLOATBUF0[24].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[25].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[25].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[25].__cell__  (.EN(\BYTE[3].FLOATBUF0[25].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[26].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[26].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[26].__cell__  (.EN(\BYTE[3].FLOATBUF0[26].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[27].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[27].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[27].__cell__  (.EN(\BYTE[3].FLOATBUF0[27].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[28].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[28].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[28].__cell__  (.EN(\BYTE[3].FLOATBUF0[28].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[29].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[29].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[29].__cell__  (.EN(\BYTE[3].FLOATBUF0[29].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[30].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[30].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[30].__cell__  (.EN(\BYTE[3].FLOATBUF0[30].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[31].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[31].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[31].__cell__  (.EN(\BYTE[3].FLOATBUF0[31].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[24].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[24].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[24].__cell__  (.EN(\BYTE[3].FLOATBUF1[24].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[25].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[25].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[25].__cell__  (.EN(\BYTE[3].FLOATBUF1[25].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[26].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[26].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[26].__cell__  (.EN(\BYTE[3].FLOATBUF1[26].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[27].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[27].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[27].__cell__  (.EN(\BYTE[3].FLOATBUF1[27].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[28].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[28].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[28].__cell__  (.EN(\BYTE[3].FLOATBUF1[28].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[29].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[29].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[29].__cell__  (.EN(\BYTE[3].FLOATBUF1[29].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[30].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[30].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[30].__cell__  (.EN(\BYTE[3].FLOATBUF1[30].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[31].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[31].TE_BN ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[31].__cell__  (.EN(\BYTE[3].FLOATBUF1[31].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \CLKBUF.__cell__  (.I(CLK),
    .Z(\CLKBUF.X ));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 \DEC0.AND0  (.A1(\A0BUF[3].X ),
    .A2(\A0BUF[4].X ),
    .A3(\DEC0.EN_N ),
    .ZN(\SLICE[0].RAM8.DEC0.EN ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC0.AND1  (.A1(\DEC0.A_N[1] ),
    .A2(\A0BUF[3].X ),
    .A3(\DEC0.EN ),
    .Z(\SLICE[1].RAM8.DEC0.EN ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC0.AND2  (.A1(\DEC0.A_N[0] ),
    .A2(\A0BUF[4].X ),
    .A3(\DEC0.EN ),
    .Z(\SLICE[2].RAM8.DEC0.EN ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC0.AND3  (.A1(\A0BUF[4].X ),
    .A2(\A0BUF[3].X ),
    .A3(\DEC0.EN ),
    .Z(\SLICE[3].RAM8.DEC0.EN ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC0.INV1  (.I(\A0BUF[3].X ),
    .ZN(\DEC0.A_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC0.INV2  (.I(\A0BUF[4].X ),
    .ZN(\DEC0.A_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC0.INV3  (.I(\DEC0.EN ),
    .ZN(\DEC0.EN_N ));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 \DEC1.AND0  (.A1(\A1BUF[3].X ),
    .A2(\A1BUF[4].X ),
    .A3(\DEC1.EN_N ),
    .ZN(\SLICE[0].RAM8.DEC1.EN ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC1.AND1  (.A1(\DEC1.A_N[1] ),
    .A2(\A1BUF[3].X ),
    .A3(\DEC1.EN ),
    .Z(\SLICE[1].RAM8.DEC1.EN ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC1.AND2  (.A1(\DEC1.A_N[0] ),
    .A2(\A1BUF[4].X ),
    .A3(\DEC1.EN ),
    .Z(\SLICE[2].RAM8.DEC1.EN ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC1.AND3  (.A1(\A1BUF[4].X ),
    .A2(\A1BUF[3].X ),
    .A3(\DEC1.EN ),
    .Z(\SLICE[3].RAM8.DEC1.EN ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC1.INV1  (.I(\A1BUF[3].X ),
    .ZN(\DEC1.A_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC1.INV2  (.I(\A1BUF[4].X ),
    .ZN(\DEC1.A_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC1.INV3  (.I(\DEC1.EN ),
    .ZN(\DEC1.EN_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[0].__cell__  (.I(Di0[0]),
    .Z(\DIBUF[0].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[10].__cell__  (.I(Di0[10]),
    .Z(\DIBUF[10].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[11].__cell__  (.I(Di0[11]),
    .Z(\DIBUF[11].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[12].__cell__  (.I(Di0[12]),
    .Z(\DIBUF[12].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[13].__cell__  (.I(Di0[13]),
    .Z(\DIBUF[13].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[14].__cell__  (.I(Di0[14]),
    .Z(\DIBUF[14].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[15].__cell__  (.I(Di0[15]),
    .Z(\DIBUF[15].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[16].__cell__  (.I(Di0[16]),
    .Z(\DIBUF[16].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[17].__cell__  (.I(Di0[17]),
    .Z(\DIBUF[17].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[18].__cell__  (.I(Di0[18]),
    .Z(\DIBUF[18].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[19].__cell__  (.I(Di0[19]),
    .Z(\DIBUF[19].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[1].__cell__  (.I(Di0[1]),
    .Z(\DIBUF[1].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[20].__cell__  (.I(Di0[20]),
    .Z(\DIBUF[20].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[21].__cell__  (.I(Di0[21]),
    .Z(\DIBUF[21].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[22].__cell__  (.I(Di0[22]),
    .Z(\DIBUF[22].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[23].__cell__  (.I(Di0[23]),
    .Z(\DIBUF[23].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[24].__cell__  (.I(Di0[24]),
    .Z(\DIBUF[24].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[25].__cell__  (.I(Di0[25]),
    .Z(\DIBUF[25].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[26].__cell__  (.I(Di0[26]),
    .Z(\DIBUF[26].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[27].__cell__  (.I(Di0[27]),
    .Z(\DIBUF[27].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[28].__cell__  (.I(Di0[28]),
    .Z(\DIBUF[28].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[29].__cell__  (.I(Di0[29]),
    .Z(\DIBUF[29].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[2].__cell__  (.I(Di0[2]),
    .Z(\DIBUF[2].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[30].__cell__  (.I(Di0[30]),
    .Z(\DIBUF[30].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[31].__cell__  (.I(Di0[31]),
    .Z(\DIBUF[31].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[3].__cell__  (.I(Di0[3]),
    .Z(\DIBUF[3].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[4].__cell__  (.I(Di0[4]),
    .Z(\DIBUF[4].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[5].__cell__  (.I(Di0[5]),
    .Z(\DIBUF[5].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[6].__cell__  (.I(Di0[6]),
    .Z(\DIBUF[6].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[7].__cell__  (.I(Di0[7]),
    .Z(\DIBUF[7].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[8].__cell__  (.I(Di0[8]),
    .Z(\DIBUF[8].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[9].__cell__  (.I(Di0[9]),
    .Z(\DIBUF[9].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Do_CLKBUF[0]  (.I(\Do0_REG.CLK_buf ),
    .Z(\Do0_REG.CLKBUF[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Do_CLKBUF[1]  (.I(\Do0_REG.CLK_buf ),
    .Z(\Do0_REG.CLKBUF[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Do_CLKBUF[2]  (.I(\Do0_REG.CLK_buf ),
    .Z(\Do0_REG.CLKBUF[2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Do_CLKBUF[3]  (.I(\Do0_REG.CLK_buf ),
    .Z(\Do0_REG.CLKBUF[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.I(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.I(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.I(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.I(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.I(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.I(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.I(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.I(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.D(\BYTE[0].FLOATBUF0[0].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.D(\BYTE[0].FLOATBUF0[1].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.D(\BYTE[0].FLOATBUF0[2].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.D(\BYTE[0].FLOATBUF0[3].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.D(\BYTE[0].FLOATBUF0[4].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.D(\BYTE[0].FLOATBUF0[5].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.D(\BYTE[0].FLOATBUF0[6].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[6]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.D(\BYTE[0].FLOATBUF0[7].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.I(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.I(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.I(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.I(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.I(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.I(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.I(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.I(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.D(\BYTE[1].FLOATBUF0[8].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[8]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.D(\BYTE[1].FLOATBUF0[9].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[9]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.D(\BYTE[1].FLOATBUF0[10].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[10]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.D(\BYTE[1].FLOATBUF0[11].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[11]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.D(\BYTE[1].FLOATBUF0[12].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[12]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.D(\BYTE[1].FLOATBUF0[13].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[13]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.D(\BYTE[1].FLOATBUF0[14].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[14]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.D(\BYTE[1].FLOATBUF0[15].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.I(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.I(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.I(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.I(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.I(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.I(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.I(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.I(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.D(\BYTE[2].FLOATBUF0[16].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[16]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.D(\BYTE[2].FLOATBUF0[17].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[17]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.D(\BYTE[2].FLOATBUF0[18].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[18]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.D(\BYTE[2].FLOATBUF0[19].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[19]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.D(\BYTE[2].FLOATBUF0[20].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[20]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.D(\BYTE[2].FLOATBUF0[21].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[21]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.D(\BYTE[2].FLOATBUF0[22].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[22]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.D(\BYTE[2].FLOATBUF0[23].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.I(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.I(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.I(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.I(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.I(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.I(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.I(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.I(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.D(\BYTE[3].FLOATBUF0[24].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[24]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.D(\BYTE[3].FLOATBUF0[25].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[25]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.D(\BYTE[3].FLOATBUF0[26].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[26]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.D(\BYTE[3].FLOATBUF0[27].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[27]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.D(\BYTE[3].FLOATBUF0[28].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[28]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.D(\BYTE[3].FLOATBUF0[29].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[29]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.D(\BYTE[3].FLOATBUF0[30].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[30]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.D(\BYTE[3].FLOATBUF0[31].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Root_CLKBUF  (.I(\CLKBUF.X ),
    .Z(\Do0_REG.CLK_buf ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Do_CLKBUF[0]  (.I(\Do1_REG.CLK_buf ),
    .Z(\Do1_REG.CLKBUF[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Do_CLKBUF[1]  (.I(\Do1_REG.CLK_buf ),
    .Z(\Do1_REG.CLKBUF[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Do_CLKBUF[2]  (.I(\Do1_REG.CLK_buf ),
    .Z(\Do1_REG.CLKBUF[2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Do_CLKBUF[3]  (.I(\Do1_REG.CLK_buf ),
    .Z(\Do1_REG.CLKBUF[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[0]  (.I(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[1]  (.I(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[2]  (.I(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[3]  (.I(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[4]  (.I(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[5]  (.I(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[6]  (.I(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[7]  (.I(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[0]  (.D(\BYTE[0].FLOATBUF1[0].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[1]  (.D(\BYTE[0].FLOATBUF1[1].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[2]  (.D(\BYTE[0].FLOATBUF1[2].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[3]  (.D(\BYTE[0].FLOATBUF1[3].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[4]  (.D(\BYTE[0].FLOATBUF1[4].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[5]  (.D(\BYTE[0].FLOATBUF1[5].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[6]  (.D(\BYTE[0].FLOATBUF1[6].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[6]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[7]  (.D(\BYTE[0].FLOATBUF1[7].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[0]  (.I(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[1]  (.I(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[2]  (.I(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[3]  (.I(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[4]  (.I(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[5]  (.I(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[6]  (.I(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[7]  (.I(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[0]  (.D(\BYTE[1].FLOATBUF1[8].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[8]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[1]  (.D(\BYTE[1].FLOATBUF1[9].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[9]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[2]  (.D(\BYTE[1].FLOATBUF1[10].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[10]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[3]  (.D(\BYTE[1].FLOATBUF1[11].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[11]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[4]  (.D(\BYTE[1].FLOATBUF1[12].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[12]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[5]  (.D(\BYTE[1].FLOATBUF1[13].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[13]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[6]  (.D(\BYTE[1].FLOATBUF1[14].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[14]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[7]  (.D(\BYTE[1].FLOATBUF1[15].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[0]  (.I(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[1]  (.I(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[2]  (.I(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[3]  (.I(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[4]  (.I(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[5]  (.I(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[6]  (.I(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[7]  (.I(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[0]  (.D(\BYTE[2].FLOATBUF1[16].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[16]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[1]  (.D(\BYTE[2].FLOATBUF1[17].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[17]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[2]  (.D(\BYTE[2].FLOATBUF1[18].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[18]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[3]  (.D(\BYTE[2].FLOATBUF1[19].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[19]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[4]  (.D(\BYTE[2].FLOATBUF1[20].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[20]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[5]  (.D(\BYTE[2].FLOATBUF1[21].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[21]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[6]  (.D(\BYTE[2].FLOATBUF1[22].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[22]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[7]  (.D(\BYTE[2].FLOATBUF1[23].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[0]  (.I(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[1]  (.I(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[2]  (.I(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[3]  (.I(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[4]  (.I(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[5]  (.I(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[6]  (.I(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[7]  (.I(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[0]  (.D(\BYTE[3].FLOATBUF1[24].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[24]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[1]  (.D(\BYTE[3].FLOATBUF1[25].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[25]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[2]  (.D(\BYTE[3].FLOATBUF1[26].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[26]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[3]  (.D(\BYTE[3].FLOATBUF1[27].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[27]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[4]  (.D(\BYTE[3].FLOATBUF1[28].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[28]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[5]  (.D(\BYTE[3].FLOATBUF1[29].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[29]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[6]  (.D(\BYTE[3].FLOATBUF1[30].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[30]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[7]  (.D(\BYTE[3].FLOATBUF1[31].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Root_CLKBUF  (.I(\CLKBUF.X ),
    .Z(\Do1_REG.CLK_buf ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \EN0BUF.__cell__  (.I(EN0),
    .Z(\DEC0.EN ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \EN1BUF.__cell__  (.I(EN1),
    .Z(\DEC1.EN ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF0[0].__cell__  (.I(EN0),
    .Z(\BYTE[0].FLOATBUF0[0].TE_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF0[1].__cell__  (.I(EN0),
    .Z(\BYTE[1].FLOATBUF0[10].TE_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF0[2].__cell__  (.I(EN0),
    .Z(\BYTE[2].FLOATBUF0[16].TE_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF0[3].__cell__  (.I(EN0),
    .Z(\BYTE[3].FLOATBUF0[24].TE_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF1[0].__cell__  (.I(EN1),
    .Z(\BYTE[0].FLOATBUF1[0].TE_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF1[1].__cell__  (.I(EN1),
    .Z(\BYTE[1].FLOATBUF1[10].TE_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF1[2].__cell__  (.I(EN1),
    .Z(\BYTE[2].FLOATBUF1[16].TE_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF1[3].__cell__  (.I(EN1),
    .Z(\BYTE[3].FLOATBUF1[24].TE_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.CLKBUF.__cell__  (.I(\CLKBUF.X ),
    .Z(\SLICE[0].RAM8.CLKBUF.X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[0]  (.I(\A0BUF[0].X ),
    .Z(\SLICE[0].RAM8.DEC0.A_buf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[1]  (.I(\A0BUF[1].X ),
    .Z(\SLICE[0].RAM8.DEC0.A_buf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[2]  (.I(\A0BUF[2].X ),
    .Z(\SLICE[0].RAM8.DEC0.A_buf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[0].RAM8.DEC0.AND0  (.A1(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf_N ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND1  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[1].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND2  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC0.A_buf_N[0] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[2].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND3  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[3].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND4  (.A1(\SLICE[0].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[4].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND5  (.A1(\SLICE[0].RAM8.DEC0.A_buf_N[1] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[5].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND6  (.A1(\SLICE[0].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[6].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND7  (.A1(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[7].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC0.ENBUF  (.I(\SLICE[0].RAM8.DEC0.EN ),
    .Z(\SLICE[0].RAM8.DEC0.EN_buf ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC0.INV1  (.I(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .ZN(\SLICE[0].RAM8.DEC0.A_buf_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC0.INV2  (.I(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[0].RAM8.DEC0.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC0.INV3  (.I(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[0].RAM8.DEC0.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC0.INV4  (.I(\SLICE[0].RAM8.DEC0.EN_buf ),
    .ZN(\SLICE[0].RAM8.DEC0.EN_buf_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[0]  (.I(\A1BUF[0].X ),
    .Z(\SLICE[0].RAM8.DEC1.A_buf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[1]  (.I(\A1BUF[1].X ),
    .Z(\SLICE[0].RAM8.DEC1.A_buf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[2]  (.I(\A1BUF[2].X ),
    .Z(\SLICE[0].RAM8.DEC1.A_buf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[0].RAM8.DEC1.AND0  (.A1(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf_N ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND1  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[1].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND2  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC1.A_buf_N[0] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[2].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND3  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[3].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND4  (.A1(\SLICE[0].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[4].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND5  (.A1(\SLICE[0].RAM8.DEC1.A_buf_N[1] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[5].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND6  (.A1(\SLICE[0].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[6].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND7  (.A1(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[7].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC1.ENBUF  (.I(\SLICE[0].RAM8.DEC1.EN ),
    .Z(\SLICE[0].RAM8.DEC1.EN_buf ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC1.INV1  (.I(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .ZN(\SLICE[0].RAM8.DEC1.A_buf_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC1.INV2  (.I(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[0].RAM8.DEC1.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC1.INV3  (.I(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[0].RAM8.DEC1.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC1.INV4  (.I(\SLICE[0].RAM8.DEC1.EN_buf ),
    .ZN(\SLICE[0].RAM8.DEC1.EN_buf_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WEBUF[0].__cell__  (.I(\SLICE[0].RAM8.WEBUF[0].A ),
    .Z(\SLICE[0].RAM8.WEBUF[0].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WEBUF[1].__cell__  (.I(\SLICE[0].RAM8.WEBUF[1].A ),
    .Z(\SLICE[0].RAM8.WEBUF[1].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WEBUF[2].__cell__  (.I(\SLICE[0].RAM8.WEBUF[2].A ),
    .Z(\SLICE[0].RAM8.WEBUF[2].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WEBUF[3].__cell__  (.I(\SLICE[0].RAM8.WEBUF[3].A ),
    .Z(\SLICE[0].RAM8.WEBUF[3].X ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[0].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[0].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[0].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[1].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[1].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[1].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[2].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[2].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[2].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[3].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[3].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[3].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[4].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[4].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[4].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[5].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[5].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[5].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[6].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[6].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[6].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[7].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[7].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[7].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.CLKBUF.__cell__  (.I(\CLKBUF.X ),
    .Z(\SLICE[1].RAM8.CLKBUF.X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[0]  (.I(\A0BUF[0].X ),
    .Z(\SLICE[1].RAM8.DEC0.A_buf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[1]  (.I(\A0BUF[1].X ),
    .Z(\SLICE[1].RAM8.DEC0.A_buf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[2]  (.I(\A0BUF[2].X ),
    .Z(\SLICE[1].RAM8.DEC0.A_buf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[1].RAM8.DEC0.AND0  (.A1(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf_N ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND1  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[1].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND2  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC0.A_buf_N[0] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[2].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND3  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[3].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND4  (.A1(\SLICE[1].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[4].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND5  (.A1(\SLICE[1].RAM8.DEC0.A_buf_N[1] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[5].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND6  (.A1(\SLICE[1].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[6].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND7  (.A1(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[7].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC0.ENBUF  (.I(\SLICE[1].RAM8.DEC0.EN ),
    .Z(\SLICE[1].RAM8.DEC0.EN_buf ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC0.INV1  (.I(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .ZN(\SLICE[1].RAM8.DEC0.A_buf_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC0.INV2  (.I(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[1].RAM8.DEC0.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC0.INV3  (.I(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[1].RAM8.DEC0.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC0.INV4  (.I(\SLICE[1].RAM8.DEC0.EN_buf ),
    .ZN(\SLICE[1].RAM8.DEC0.EN_buf_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[0]  (.I(\A1BUF[0].X ),
    .Z(\SLICE[1].RAM8.DEC1.A_buf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[1]  (.I(\A1BUF[1].X ),
    .Z(\SLICE[1].RAM8.DEC1.A_buf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[2]  (.I(\A1BUF[2].X ),
    .Z(\SLICE[1].RAM8.DEC1.A_buf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[1].RAM8.DEC1.AND0  (.A1(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf_N ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND1  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[1].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND2  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC1.A_buf_N[0] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[2].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND3  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[3].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND4  (.A1(\SLICE[1].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[4].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND5  (.A1(\SLICE[1].RAM8.DEC1.A_buf_N[1] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[5].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND6  (.A1(\SLICE[1].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[6].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND7  (.A1(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[7].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC1.ENBUF  (.I(\SLICE[1].RAM8.DEC1.EN ),
    .Z(\SLICE[1].RAM8.DEC1.EN_buf ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC1.INV1  (.I(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .ZN(\SLICE[1].RAM8.DEC1.A_buf_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC1.INV2  (.I(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[1].RAM8.DEC1.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC1.INV3  (.I(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[1].RAM8.DEC1.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC1.INV4  (.I(\SLICE[1].RAM8.DEC1.EN_buf ),
    .ZN(\SLICE[1].RAM8.DEC1.EN_buf_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WEBUF[0].__cell__  (.I(\SLICE[0].RAM8.WEBUF[0].A ),
    .Z(\SLICE[1].RAM8.WEBUF[0].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WEBUF[1].__cell__  (.I(\SLICE[0].RAM8.WEBUF[1].A ),
    .Z(\SLICE[1].RAM8.WEBUF[1].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WEBUF[2].__cell__  (.I(\SLICE[0].RAM8.WEBUF[2].A ),
    .Z(\SLICE[1].RAM8.WEBUF[2].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WEBUF[3].__cell__  (.I(\SLICE[0].RAM8.WEBUF[3].A ),
    .Z(\SLICE[1].RAM8.WEBUF[3].X ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[0].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[0].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[0].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[1].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[1].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[1].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[2].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[2].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[2].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[3].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[3].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[3].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[4].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[4].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[4].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[5].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[5].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[5].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[6].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[6].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[6].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[7].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[7].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[7].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.CLKBUF.__cell__  (.I(\CLKBUF.X ),
    .Z(\SLICE[2].RAM8.CLKBUF.X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[0]  (.I(\A0BUF[0].X ),
    .Z(\SLICE[2].RAM8.DEC0.A_buf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[1]  (.I(\A0BUF[1].X ),
    .Z(\SLICE[2].RAM8.DEC0.A_buf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[2]  (.I(\A0BUF[2].X ),
    .Z(\SLICE[2].RAM8.DEC0.A_buf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[2].RAM8.DEC0.AND0  (.A1(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf_N ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND1  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[1].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND2  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC0.A_buf_N[0] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[2].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND3  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[3].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND4  (.A1(\SLICE[2].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[4].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND5  (.A1(\SLICE[2].RAM8.DEC0.A_buf_N[1] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[5].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND6  (.A1(\SLICE[2].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[6].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND7  (.A1(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[7].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC0.ENBUF  (.I(\SLICE[2].RAM8.DEC0.EN ),
    .Z(\SLICE[2].RAM8.DEC0.EN_buf ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC0.INV1  (.I(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .ZN(\SLICE[2].RAM8.DEC0.A_buf_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC0.INV2  (.I(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[2].RAM8.DEC0.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC0.INV3  (.I(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[2].RAM8.DEC0.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC0.INV4  (.I(\SLICE[2].RAM8.DEC0.EN_buf ),
    .ZN(\SLICE[2].RAM8.DEC0.EN_buf_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[0]  (.I(\A1BUF[0].X ),
    .Z(\SLICE[2].RAM8.DEC1.A_buf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[1]  (.I(\A1BUF[1].X ),
    .Z(\SLICE[2].RAM8.DEC1.A_buf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[2]  (.I(\A1BUF[2].X ),
    .Z(\SLICE[2].RAM8.DEC1.A_buf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[2].RAM8.DEC1.AND0  (.A1(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf_N ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND1  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[1].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND2  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC1.A_buf_N[0] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[2].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND3  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[3].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND4  (.A1(\SLICE[2].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[4].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND5  (.A1(\SLICE[2].RAM8.DEC1.A_buf_N[1] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[5].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND6  (.A1(\SLICE[2].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[6].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND7  (.A1(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[7].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC1.ENBUF  (.I(\SLICE[2].RAM8.DEC1.EN ),
    .Z(\SLICE[2].RAM8.DEC1.EN_buf ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC1.INV1  (.I(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .ZN(\SLICE[2].RAM8.DEC1.A_buf_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC1.INV2  (.I(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[2].RAM8.DEC1.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC1.INV3  (.I(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[2].RAM8.DEC1.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC1.INV4  (.I(\SLICE[2].RAM8.DEC1.EN_buf ),
    .ZN(\SLICE[2].RAM8.DEC1.EN_buf_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WEBUF[0].__cell__  (.I(\SLICE[0].RAM8.WEBUF[0].A ),
    .Z(\SLICE[2].RAM8.WEBUF[0].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WEBUF[1].__cell__  (.I(\SLICE[0].RAM8.WEBUF[1].A ),
    .Z(\SLICE[2].RAM8.WEBUF[1].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WEBUF[2].__cell__  (.I(\SLICE[0].RAM8.WEBUF[2].A ),
    .Z(\SLICE[2].RAM8.WEBUF[2].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WEBUF[3].__cell__  (.I(\SLICE[0].RAM8.WEBUF[3].A ),
    .Z(\SLICE[2].RAM8.WEBUF[3].X ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[0].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[0].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[0].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[0].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[0].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[1].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[1].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[1].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[1].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[1].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[2].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[2].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[2].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[2].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[2].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[3].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[3].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[3].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[3].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[3].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[4].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[4].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[4].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[4].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[4].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[5].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[5].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[5].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[5].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[5].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[6].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[6].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[6].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[6].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[6].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[7].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[7].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[7].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[7].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[7].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.CLKBUF.__cell__  (.I(\CLKBUF.X ),
    .Z(\SLICE[3].RAM8.CLKBUF.X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[0]  (.I(\A0BUF[0].X ),
    .Z(\SLICE[3].RAM8.DEC0.A_buf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[1]  (.I(\A0BUF[1].X ),
    .Z(\SLICE[3].RAM8.DEC0.A_buf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[2]  (.I(\A0BUF[2].X ),
    .Z(\SLICE[3].RAM8.DEC0.A_buf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[3].RAM8.DEC0.AND0  (.A1(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf_N ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND1  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[1].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND2  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC0.A_buf_N[0] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[2].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND3  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[3].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND4  (.A1(\SLICE[3].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[4].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND5  (.A1(\SLICE[3].RAM8.DEC0.A_buf_N[1] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[5].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND6  (.A1(\SLICE[3].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[6].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND7  (.A1(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[7].W.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC0.ENBUF  (.I(\SLICE[3].RAM8.DEC0.EN ),
    .Z(\SLICE[3].RAM8.DEC0.EN_buf ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC0.INV1  (.I(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .ZN(\SLICE[3].RAM8.DEC0.A_buf_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC0.INV2  (.I(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[3].RAM8.DEC0.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC0.INV3  (.I(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[3].RAM8.DEC0.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC0.INV4  (.I(\SLICE[3].RAM8.DEC0.EN_buf ),
    .ZN(\SLICE[3].RAM8.DEC0.EN_buf_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[0]  (.I(\A1BUF[0].X ),
    .Z(\SLICE[3].RAM8.DEC1.A_buf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[1]  (.I(\A1BUF[1].X ),
    .Z(\SLICE[3].RAM8.DEC1.A_buf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[2]  (.I(\A1BUF[2].X ),
    .Z(\SLICE[3].RAM8.DEC1.A_buf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[3].RAM8.DEC1.AND0  (.A1(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf_N ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND1  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[1].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND2  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC1.A_buf_N[0] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[2].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND3  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[3].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND4  (.A1(\SLICE[3].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[4].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND5  (.A1(\SLICE[3].RAM8.DEC1.A_buf_N[1] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[5].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND6  (.A1(\SLICE[3].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[6].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND7  (.A1(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[7].W.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC1.ENBUF  (.I(\SLICE[3].RAM8.DEC1.EN ),
    .Z(\SLICE[3].RAM8.DEC1.EN_buf ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC1.INV1  (.I(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .ZN(\SLICE[3].RAM8.DEC1.A_buf_N[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC1.INV2  (.I(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[3].RAM8.DEC1.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC1.INV3  (.I(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[3].RAM8.DEC1.A_buf_N[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC1.INV4  (.I(\SLICE[3].RAM8.DEC1.EN_buf ),
    .ZN(\SLICE[3].RAM8.DEC1.EN_buf_N ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WEBUF[0].__cell__  (.I(\SLICE[0].RAM8.WEBUF[0].A ),
    .Z(\SLICE[3].RAM8.WEBUF[0].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WEBUF[1].__cell__  (.I(\SLICE[0].RAM8.WEBUF[1].A ),
    .Z(\SLICE[3].RAM8.WEBUF[1].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WEBUF[2].__cell__  (.I(\SLICE[0].RAM8.WEBUF[2].A ),
    .Z(\SLICE[3].RAM8.WEBUF[2].X ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WEBUF[3].__cell__  (.I(\SLICE[0].RAM8.WEBUF[3].A ),
    .Z(\SLICE[3].RAM8.WEBUF[3].X ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[0].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[0].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[0].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[0].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[0].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[1].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[1].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[1].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[1].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[1].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[2].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[2].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[2].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[2].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[2].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[3].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[3].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[3].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[3].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[3].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[4].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[4].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[4].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[4].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[4].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[5].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[5].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[5].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[5].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[5].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[6].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[6].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[6].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[6].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[6].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[7].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[7].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[7].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[7].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[7].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE0[0].__cell__  (.ZN(\BYTE[0].FLOATBUF0[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE0[1].__cell__  (.ZN(\BYTE[1].FLOATBUF0[10].A ));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE0[2].__cell__  (.ZN(\BYTE[2].FLOATBUF0[16].A ));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE0[3].__cell__  (.ZN(\BYTE[3].FLOATBUF0[24].A ));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE1[0].__cell__  (.ZN(\BYTE[0].FLOATBUF1[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE1[1].__cell__  (.ZN(\BYTE[1].FLOATBUF1[10].A ));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE1[2].__cell__  (.ZN(\BYTE[2].FLOATBUF1[16].A ));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE1[3].__cell__  (.ZN(\BYTE[3].FLOATBUF1[24].A ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \WEBUF[0].__cell__  (.I(WE0[0]),
    .Z(\SLICE[0].RAM8.WEBUF[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \WEBUF[1].__cell__  (.I(WE0[1]),
    .Z(\SLICE[0].RAM8.WEBUF[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \WEBUF[2].__cell__  (.I(WE0[2]),
    .Z(\SLICE[0].RAM8.WEBUF[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \WEBUF[3].__cell__  (.I(WE0[3]),
    .Z(\SLICE[0].RAM8.WEBUF[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__tiel TIE_ZERO_zero_ (.ZN(zero_));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_0_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_1_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_2_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_3_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_4_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_5_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_8_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_10_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_11_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_12_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_13_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_14_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_15_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_16_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_2_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_3_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_4_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_5_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_5_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_6_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_7_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_8_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_8_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_6_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_7_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_10_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_10_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_11_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_12_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_12_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_13_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_13_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_14_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_14_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_15_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_15_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_16_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_16_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_14_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_15_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_16_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_18_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_19_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_20_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_21_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_22_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_23_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_24_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_22_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_23_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_24_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_26_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_27_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_28_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_29_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_30_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_31_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_32_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_30_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_31_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_32_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_0 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_1 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_3 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_4 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_5 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_0_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_0_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_0_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_1_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_2_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_2_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_2_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_2_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_2_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_3_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_3_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_3_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_3_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_4_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_4_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_4_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_4_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_4_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_5_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_5_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_5_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_5_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_5_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_6_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_6_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_6_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_6_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_7_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_7_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_7_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_7_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_8_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_8_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_8_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_8_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_8_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_9_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_9_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_9_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_9_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_9_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_10_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_10_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_10_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_11_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_11_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_11_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_11_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_12_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_12_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_12_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_12_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_12_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_13_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_13_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_13_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_13_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_13_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_14_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_14_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_14_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_14_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_15_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_15_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_15_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_16_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_16_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_16_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_16_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_17_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_17_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_18_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_18_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_18_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_18_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_19_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_19_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_19_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_19_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_20_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_20_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_20_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_21_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_21_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_21_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_21_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_22_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_22_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_22_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_23_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_23_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_23_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_23_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_23_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_24_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_24_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_24_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_24_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_25_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_25_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_25_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_25_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_25_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_26_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_26_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_26_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_26_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_27_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_27_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_27_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_28_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_28_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_28_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_28_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_28_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_29_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_29_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_29_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_29_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_29_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_30_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_30_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_30_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_31_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_31_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_31_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_31_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_31_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_32_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_32_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_32_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_32_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_0 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_1 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_3 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_33_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_33_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_33_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_33_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_33_802 ();
endmodule

