magic
tech gf180mcuC
magscale 1 5
timestamp 1676188205
<< obsm1 >>
rect 233 15 127176 16057
<< metal2 >>
rect 1960 15872 2016 16072
rect 3920 15872 3976 16072
rect 5880 15872 5936 16072
rect 7840 15872 7896 16072
rect 9800 15872 9856 16072
rect 11760 15872 11816 16072
rect 13720 15872 13776 16072
rect 15680 15872 15736 16072
rect 17640 15872 17696 16072
rect 19600 15872 19656 16072
rect 21560 15872 21616 16072
rect 23520 15872 23576 16072
rect 25480 15872 25536 16072
rect 27440 15872 27496 16072
rect 29400 15872 29456 16072
rect 31360 15872 31416 16072
rect 33320 15872 33376 16072
rect 35280 15872 35336 16072
rect 37240 15872 37296 16072
rect 39200 15872 39256 16072
rect 41160 15872 41216 16072
rect 43120 15872 43176 16072
rect 45080 15872 45136 16072
rect 47040 15872 47096 16072
rect 49000 15872 49056 16072
rect 50960 15872 51016 16072
rect 52920 15872 52976 16072
rect 54880 15872 54936 16072
rect 56840 15872 56896 16072
rect 58800 15872 58856 16072
rect 60760 15872 60816 16072
rect 62720 15872 62776 16072
rect 64680 15872 64736 16072
rect 66640 15872 66696 16072
rect 68600 15872 68656 16072
rect 70560 15872 70616 16072
rect 72520 15872 72576 16072
rect 74480 15872 74536 16072
rect 76440 15872 76496 16072
rect 78400 15872 78456 16072
rect 80360 15872 80416 16072
rect 82320 15872 82376 16072
rect 84280 15872 84336 16072
rect 86240 15872 86296 16072
rect 88200 15872 88256 16072
rect 90160 15872 90216 16072
rect 92120 15872 92176 16072
rect 94080 15872 94136 16072
rect 96040 15872 96096 16072
rect 98000 15872 98056 16072
rect 99960 15872 100016 16072
rect 101920 15872 101976 16072
rect 103880 15872 103936 16072
rect 105840 15872 105896 16072
rect 107800 15872 107856 16072
rect 109760 15872 109816 16072
rect 111720 15872 111776 16072
rect 113680 15872 113736 16072
rect 115640 15872 115696 16072
rect 117600 15872 117656 16072
rect 119560 15872 119616 16072
rect 121520 15872 121576 16072
rect 123480 15872 123536 16072
rect 125440 15872 125496 16072
rect 2072 0 2128 200
rect 6048 0 6104 200
rect 10024 0 10080 200
rect 14000 0 14056 200
rect 17976 0 18032 200
rect 21952 0 22008 200
rect 25928 0 25984 200
rect 29904 0 29960 200
rect 33880 0 33936 200
rect 37856 0 37912 200
rect 41832 0 41888 200
rect 45808 0 45864 200
rect 49784 0 49840 200
rect 53760 0 53816 200
rect 57736 0 57792 200
rect 61712 0 61768 200
rect 65688 0 65744 200
rect 69664 0 69720 200
rect 73640 0 73696 200
rect 77616 0 77672 200
rect 81592 0 81648 200
rect 85568 0 85624 200
rect 89544 0 89600 200
rect 93520 0 93576 200
rect 97496 0 97552 200
rect 101472 0 101528 200
rect 105448 0 105504 200
rect 109424 0 109480 200
rect 113400 0 113456 200
rect 117376 0 117432 200
rect 121352 0 121408 200
rect 125328 0 125384 200
<< obsm2 >>
rect 14 15842 1930 16063
rect 2046 15842 3890 16063
rect 4006 15842 5850 16063
rect 5966 15842 7810 16063
rect 7926 15842 9770 16063
rect 9886 15842 11730 16063
rect 11846 15842 13690 16063
rect 13806 15842 15650 16063
rect 15766 15842 17610 16063
rect 17726 15842 19570 16063
rect 19686 15842 21530 16063
rect 21646 15842 23490 16063
rect 23606 15842 25450 16063
rect 25566 15842 27410 16063
rect 27526 15842 29370 16063
rect 29486 15842 31330 16063
rect 31446 15842 33290 16063
rect 33406 15842 35250 16063
rect 35366 15842 37210 16063
rect 37326 15842 39170 16063
rect 39286 15842 41130 16063
rect 41246 15842 43090 16063
rect 43206 15842 45050 16063
rect 45166 15842 47010 16063
rect 47126 15842 48970 16063
rect 49086 15842 50930 16063
rect 51046 15842 52890 16063
rect 53006 15842 54850 16063
rect 54966 15842 56810 16063
rect 56926 15842 58770 16063
rect 58886 15842 60730 16063
rect 60846 15842 62690 16063
rect 62806 15842 64650 16063
rect 64766 15842 66610 16063
rect 66726 15842 68570 16063
rect 68686 15842 70530 16063
rect 70646 15842 72490 16063
rect 72606 15842 74450 16063
rect 74566 15842 76410 16063
rect 76526 15842 78370 16063
rect 78486 15842 80330 16063
rect 80446 15842 82290 16063
rect 82406 15842 84250 16063
rect 84366 15842 86210 16063
rect 86326 15842 88170 16063
rect 88286 15842 90130 16063
rect 90246 15842 92090 16063
rect 92206 15842 94050 16063
rect 94166 15842 96010 16063
rect 96126 15842 97970 16063
rect 98086 15842 99930 16063
rect 100046 15842 101890 16063
rect 102006 15842 103850 16063
rect 103966 15842 105810 16063
rect 105926 15842 107770 16063
rect 107886 15842 109730 16063
rect 109846 15842 111690 16063
rect 111806 15842 113650 16063
rect 113766 15842 115610 16063
rect 115726 15842 117570 16063
rect 117686 15842 119530 16063
rect 119646 15842 121490 16063
rect 121606 15842 123450 16063
rect 123566 15842 125410 16063
rect 125526 15842 127330 16063
rect 14 230 127330 15842
rect 14 9 2042 230
rect 2158 9 6018 230
rect 6134 9 9994 230
rect 10110 9 13970 230
rect 14086 9 17946 230
rect 18062 9 21922 230
rect 22038 9 25898 230
rect 26014 9 29874 230
rect 29990 9 33850 230
rect 33966 9 37826 230
rect 37942 9 41802 230
rect 41918 9 45778 230
rect 45894 9 49754 230
rect 49870 9 53730 230
rect 53846 9 57706 230
rect 57822 9 61682 230
rect 61798 9 65658 230
rect 65774 9 69634 230
rect 69750 9 73610 230
rect 73726 9 77586 230
rect 77702 9 81562 230
rect 81678 9 85538 230
rect 85654 9 89514 230
rect 89630 9 93490 230
rect 93606 9 97466 230
rect 97582 9 101442 230
rect 101558 9 105418 230
rect 105534 9 109394 230
rect 109510 9 113370 230
rect 113486 9 117346 230
rect 117462 9 121322 230
rect 121438 9 125298 230
rect 125414 9 127330 230
<< metal3 >>
rect 127256 15064 127456 15120
rect 0 14896 200 14952
rect 127256 13496 127456 13552
rect 0 12600 200 12656
rect 127256 11928 127456 11984
rect 0 10304 200 10360
rect 127256 10360 127456 10416
rect 127256 8792 127456 8848
rect 0 8008 200 8064
rect 127256 7224 127456 7280
rect 0 5712 200 5768
rect 127256 5656 127456 5712
rect 127256 4088 127456 4144
rect 0 3416 200 3472
rect 127256 2520 127456 2576
rect 0 1120 200 1176
rect 127256 952 127456 1008
<< obsm3 >>
rect 177 15150 127335 16058
rect 177 15034 127226 15150
rect 177 14982 127335 15034
rect 230 14866 127335 14982
rect 177 13582 127335 14866
rect 177 13466 127226 13582
rect 177 12686 127335 13466
rect 230 12570 127335 12686
rect 177 12014 127335 12570
rect 177 11898 127226 12014
rect 177 10446 127335 11898
rect 177 10390 127226 10446
rect 230 10330 127226 10390
rect 230 10274 127335 10330
rect 177 8878 127335 10274
rect 177 8762 127226 8878
rect 177 8094 127335 8762
rect 230 7978 127335 8094
rect 177 7310 127335 7978
rect 177 7194 127226 7310
rect 177 5798 127335 7194
rect 230 5742 127335 5798
rect 230 5682 127226 5742
rect 177 5626 127226 5682
rect 177 4174 127335 5626
rect 177 4058 127226 4174
rect 177 3502 127335 4058
rect 230 3386 127335 3502
rect 177 2606 127335 3386
rect 177 2490 127226 2606
rect 177 1206 127335 2490
rect 230 1090 127335 1206
rect 177 1038 127335 1090
rect 177 922 127226 1038
rect 177 14 127335 922
<< metal4 >>
rect 1832 1146 1992 14926
rect 9512 1146 9672 14926
rect 17192 1146 17352 14926
rect 24872 1146 25032 14926
rect 32552 1146 32712 14926
rect 40232 1146 40392 14926
rect 47912 1146 48072 14926
rect 55592 1146 55752 14926
rect 63272 1146 63432 14926
rect 70952 1146 71112 14926
rect 78632 1146 78792 14926
rect 86312 1146 86472 14926
rect 93992 1146 94152 14926
rect 101672 1146 101832 14926
rect 109352 1146 109512 14926
rect 117032 1146 117192 14926
rect 124712 1146 124872 14926
<< obsm4 >>
rect 350 14956 110362 16063
rect 350 1116 1802 14956
rect 2022 1116 9482 14956
rect 9702 1116 17162 14956
rect 17382 1116 24842 14956
rect 25062 1116 32522 14956
rect 32742 1116 40202 14956
rect 40422 1116 47882 14956
rect 48102 1116 55562 14956
rect 55782 1116 63242 14956
rect 63462 1116 70922 14956
rect 71142 1116 78602 14956
rect 78822 1116 86282 14956
rect 86502 1116 93962 14956
rect 94182 1116 101642 14956
rect 101862 1116 109322 14956
rect 109542 1116 110362 14956
rect 350 9 110362 1116
<< labels >>
rlabel metal3 s 127256 8792 127456 8848 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 127256 10360 127456 10416 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 127256 11928 127456 11984 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 127256 13496 127456 13552 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 127256 15064 127456 15120 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 0 3416 200 3472 6 A1[0]
port 6 nsew signal input
rlabel metal3 s 0 5712 200 5768 6 A1[1]
port 7 nsew signal input
rlabel metal3 s 0 8008 200 8064 6 A1[2]
port 8 nsew signal input
rlabel metal3 s 0 10304 200 10360 6 A1[3]
port 9 nsew signal input
rlabel metal3 s 0 12600 200 12656 6 A1[4]
port 10 nsew signal input
rlabel metal3 s 0 1120 200 1176 6 CLK
port 11 nsew signal input
rlabel metal2 s 2072 0 2128 200 6 Di0[0]
port 12 nsew signal input
rlabel metal2 s 41832 0 41888 200 6 Di0[10]
port 13 nsew signal input
rlabel metal2 s 45808 0 45864 200 6 Di0[11]
port 14 nsew signal input
rlabel metal2 s 49784 0 49840 200 6 Di0[12]
port 15 nsew signal input
rlabel metal2 s 53760 0 53816 200 6 Di0[13]
port 16 nsew signal input
rlabel metal2 s 57736 0 57792 200 6 Di0[14]
port 17 nsew signal input
rlabel metal2 s 61712 0 61768 200 6 Di0[15]
port 18 nsew signal input
rlabel metal2 s 65688 0 65744 200 6 Di0[16]
port 19 nsew signal input
rlabel metal2 s 69664 0 69720 200 6 Di0[17]
port 20 nsew signal input
rlabel metal2 s 73640 0 73696 200 6 Di0[18]
port 21 nsew signal input
rlabel metal2 s 77616 0 77672 200 6 Di0[19]
port 22 nsew signal input
rlabel metal2 s 6048 0 6104 200 6 Di0[1]
port 23 nsew signal input
rlabel metal2 s 81592 0 81648 200 6 Di0[20]
port 24 nsew signal input
rlabel metal2 s 85568 0 85624 200 6 Di0[21]
port 25 nsew signal input
rlabel metal2 s 89544 0 89600 200 6 Di0[22]
port 26 nsew signal input
rlabel metal2 s 93520 0 93576 200 6 Di0[23]
port 27 nsew signal input
rlabel metal2 s 97496 0 97552 200 6 Di0[24]
port 28 nsew signal input
rlabel metal2 s 101472 0 101528 200 6 Di0[25]
port 29 nsew signal input
rlabel metal2 s 105448 0 105504 200 6 Di0[26]
port 30 nsew signal input
rlabel metal2 s 109424 0 109480 200 6 Di0[27]
port 31 nsew signal input
rlabel metal2 s 113400 0 113456 200 6 Di0[28]
port 32 nsew signal input
rlabel metal2 s 117376 0 117432 200 6 Di0[29]
port 33 nsew signal input
rlabel metal2 s 10024 0 10080 200 6 Di0[2]
port 34 nsew signal input
rlabel metal2 s 121352 0 121408 200 6 Di0[30]
port 35 nsew signal input
rlabel metal2 s 125328 0 125384 200 6 Di0[31]
port 36 nsew signal input
rlabel metal2 s 14000 0 14056 200 6 Di0[3]
port 37 nsew signal input
rlabel metal2 s 17976 0 18032 200 6 Di0[4]
port 38 nsew signal input
rlabel metal2 s 21952 0 22008 200 6 Di0[5]
port 39 nsew signal input
rlabel metal2 s 25928 0 25984 200 6 Di0[6]
port 40 nsew signal input
rlabel metal2 s 29904 0 29960 200 6 Di0[7]
port 41 nsew signal input
rlabel metal2 s 33880 0 33936 200 6 Di0[8]
port 42 nsew signal input
rlabel metal2 s 37856 0 37912 200 6 Di0[9]
port 43 nsew signal input
rlabel metal2 s 1960 15872 2016 16072 6 Do0[0]
port 44 nsew signal output
rlabel metal2 s 21560 15872 21616 16072 6 Do0[10]
port 45 nsew signal output
rlabel metal2 s 25480 15872 25536 16072 6 Do0[11]
port 46 nsew signal output
rlabel metal2 s 29400 15872 29456 16072 6 Do0[12]
port 47 nsew signal output
rlabel metal2 s 33320 15872 33376 16072 6 Do0[13]
port 48 nsew signal output
rlabel metal2 s 37240 15872 37296 16072 6 Do0[14]
port 49 nsew signal output
rlabel metal2 s 41160 15872 41216 16072 6 Do0[15]
port 50 nsew signal output
rlabel metal2 s 45080 15872 45136 16072 6 Do0[16]
port 51 nsew signal output
rlabel metal2 s 49000 15872 49056 16072 6 Do0[17]
port 52 nsew signal output
rlabel metal2 s 52920 15872 52976 16072 6 Do0[18]
port 53 nsew signal output
rlabel metal2 s 56840 15872 56896 16072 6 Do0[19]
port 54 nsew signal output
rlabel metal2 s 3920 15872 3976 16072 6 Do0[1]
port 55 nsew signal output
rlabel metal2 s 60760 15872 60816 16072 6 Do0[20]
port 56 nsew signal output
rlabel metal2 s 62720 15872 62776 16072 6 Do0[21]
port 57 nsew signal output
rlabel metal2 s 64680 15872 64736 16072 6 Do0[22]
port 58 nsew signal output
rlabel metal2 s 66640 15872 66696 16072 6 Do0[23]
port 59 nsew signal output
rlabel metal2 s 68600 15872 68656 16072 6 Do0[24]
port 60 nsew signal output
rlabel metal2 s 70560 15872 70616 16072 6 Do0[25]
port 61 nsew signal output
rlabel metal2 s 72520 15872 72576 16072 6 Do0[26]
port 62 nsew signal output
rlabel metal2 s 74480 15872 74536 16072 6 Do0[27]
port 63 nsew signal output
rlabel metal2 s 76440 15872 76496 16072 6 Do0[28]
port 64 nsew signal output
rlabel metal2 s 78400 15872 78456 16072 6 Do0[29]
port 65 nsew signal output
rlabel metal2 s 5880 15872 5936 16072 6 Do0[2]
port 66 nsew signal output
rlabel metal2 s 80360 15872 80416 16072 6 Do0[30]
port 67 nsew signal output
rlabel metal2 s 82320 15872 82376 16072 6 Do0[31]
port 68 nsew signal output
rlabel metal2 s 7840 15872 7896 16072 6 Do0[3]
port 69 nsew signal output
rlabel metal2 s 9800 15872 9856 16072 6 Do0[4]
port 70 nsew signal output
rlabel metal2 s 11760 15872 11816 16072 6 Do0[5]
port 71 nsew signal output
rlabel metal2 s 13720 15872 13776 16072 6 Do0[6]
port 72 nsew signal output
rlabel metal2 s 15680 15872 15736 16072 6 Do0[7]
port 73 nsew signal output
rlabel metal2 s 17640 15872 17696 16072 6 Do0[8]
port 74 nsew signal output
rlabel metal2 s 19600 15872 19656 16072 6 Do0[9]
port 75 nsew signal output
rlabel metal2 s 23520 15872 23576 16072 6 Do1[0]
port 76 nsew signal output
rlabel metal2 s 84280 15872 84336 16072 6 Do1[10]
port 77 nsew signal output
rlabel metal2 s 86240 15872 86296 16072 6 Do1[11]
port 78 nsew signal output
rlabel metal2 s 88200 15872 88256 16072 6 Do1[12]
port 79 nsew signal output
rlabel metal2 s 90160 15872 90216 16072 6 Do1[13]
port 80 nsew signal output
rlabel metal2 s 92120 15872 92176 16072 6 Do1[14]
port 81 nsew signal output
rlabel metal2 s 94080 15872 94136 16072 6 Do1[15]
port 82 nsew signal output
rlabel metal2 s 96040 15872 96096 16072 6 Do1[16]
port 83 nsew signal output
rlabel metal2 s 98000 15872 98056 16072 6 Do1[17]
port 84 nsew signal output
rlabel metal2 s 99960 15872 100016 16072 6 Do1[18]
port 85 nsew signal output
rlabel metal2 s 101920 15872 101976 16072 6 Do1[19]
port 86 nsew signal output
rlabel metal2 s 27440 15872 27496 16072 6 Do1[1]
port 87 nsew signal output
rlabel metal2 s 103880 15872 103936 16072 6 Do1[20]
port 88 nsew signal output
rlabel metal2 s 105840 15872 105896 16072 6 Do1[21]
port 89 nsew signal output
rlabel metal2 s 107800 15872 107856 16072 6 Do1[22]
port 90 nsew signal output
rlabel metal2 s 109760 15872 109816 16072 6 Do1[23]
port 91 nsew signal output
rlabel metal2 s 111720 15872 111776 16072 6 Do1[24]
port 92 nsew signal output
rlabel metal2 s 113680 15872 113736 16072 6 Do1[25]
port 93 nsew signal output
rlabel metal2 s 115640 15872 115696 16072 6 Do1[26]
port 94 nsew signal output
rlabel metal2 s 117600 15872 117656 16072 6 Do1[27]
port 95 nsew signal output
rlabel metal2 s 119560 15872 119616 16072 6 Do1[28]
port 96 nsew signal output
rlabel metal2 s 121520 15872 121576 16072 6 Do1[29]
port 97 nsew signal output
rlabel metal2 s 31360 15872 31416 16072 6 Do1[2]
port 98 nsew signal output
rlabel metal2 s 123480 15872 123536 16072 6 Do1[30]
port 99 nsew signal output
rlabel metal2 s 125440 15872 125496 16072 6 Do1[31]
port 100 nsew signal output
rlabel metal2 s 35280 15872 35336 16072 6 Do1[3]
port 101 nsew signal output
rlabel metal2 s 39200 15872 39256 16072 6 Do1[4]
port 102 nsew signal output
rlabel metal2 s 43120 15872 43176 16072 6 Do1[5]
port 103 nsew signal output
rlabel metal2 s 47040 15872 47096 16072 6 Do1[6]
port 104 nsew signal output
rlabel metal2 s 50960 15872 51016 16072 6 Do1[7]
port 105 nsew signal output
rlabel metal2 s 54880 15872 54936 16072 6 Do1[8]
port 106 nsew signal output
rlabel metal2 s 58800 15872 58856 16072 6 Do1[9]
port 107 nsew signal output
rlabel metal3 s 127256 952 127456 1008 6 EN0
port 108 nsew signal input
rlabel metal3 s 0 14896 200 14952 6 EN1
port 109 nsew signal input
rlabel metal4 s 1832 1146 1992 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 17192 1146 17352 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 32552 1146 32712 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 47912 1146 48072 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 63272 1146 63432 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 78632 1146 78792 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 93992 1146 94152 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 109352 1146 109512 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 124712 1146 124872 14926 6 VDD
port 110 nsew power bidirectional
rlabel metal4 s 9512 1146 9672 14926 6 VSS
port 111 nsew ground bidirectional
rlabel metal4 s 24872 1146 25032 14926 6 VSS
port 111 nsew ground bidirectional
rlabel metal4 s 40232 1146 40392 14926 6 VSS
port 111 nsew ground bidirectional
rlabel metal4 s 55592 1146 55752 14926 6 VSS
port 111 nsew ground bidirectional
rlabel metal4 s 70952 1146 71112 14926 6 VSS
port 111 nsew ground bidirectional
rlabel metal4 s 86312 1146 86472 14926 6 VSS
port 111 nsew ground bidirectional
rlabel metal4 s 101672 1146 101832 14926 6 VSS
port 111 nsew ground bidirectional
rlabel metal4 s 117032 1146 117192 14926 6 VSS
port 111 nsew ground bidirectional
rlabel metal3 s 127256 2520 127456 2576 6 WE0[0]
port 112 nsew signal input
rlabel metal3 s 127256 4088 127456 4144 6 WE0[1]
port 113 nsew signal input
rlabel metal3 s 127256 5656 127456 5712 6 WE0[2]
port 114 nsew signal input
rlabel metal3 s 127256 7224 127456 7280 6 WE0[3]
port 115 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 127456 16072
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8730990
string GDS_FILE /si/work/DFFRAM/build/32x32_1RW1R/openlane/runs/RUN_2023.02.12_15.34.01/results/signoff/RAM32_1RW1R.magic.gds
string GDS_START 94508
<< end >>

