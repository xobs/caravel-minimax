// This is the unpowered netlist.
module minimax_rf (clk,
    we,
    addrD,
    addrS,
    new_value,
    rD,
    rS);
 input clk;
 input we;
 input [4:0] addrD;
 input [4:0] addrS;
 input [31:0] new_value;
 output [31:0] rD;
 output [31:0] rS;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire \register_file[10][0] ;
 wire \register_file[10][10] ;
 wire \register_file[10][11] ;
 wire \register_file[10][12] ;
 wire \register_file[10][13] ;
 wire \register_file[10][14] ;
 wire \register_file[10][15] ;
 wire \register_file[10][16] ;
 wire \register_file[10][17] ;
 wire \register_file[10][18] ;
 wire \register_file[10][19] ;
 wire \register_file[10][1] ;
 wire \register_file[10][20] ;
 wire \register_file[10][21] ;
 wire \register_file[10][22] ;
 wire \register_file[10][23] ;
 wire \register_file[10][24] ;
 wire \register_file[10][25] ;
 wire \register_file[10][26] ;
 wire \register_file[10][27] ;
 wire \register_file[10][28] ;
 wire \register_file[10][29] ;
 wire \register_file[10][2] ;
 wire \register_file[10][30] ;
 wire \register_file[10][31] ;
 wire \register_file[10][3] ;
 wire \register_file[10][4] ;
 wire \register_file[10][5] ;
 wire \register_file[10][6] ;
 wire \register_file[10][7] ;
 wire \register_file[10][8] ;
 wire \register_file[10][9] ;
 wire \register_file[11][0] ;
 wire \register_file[11][10] ;
 wire \register_file[11][11] ;
 wire \register_file[11][12] ;
 wire \register_file[11][13] ;
 wire \register_file[11][14] ;
 wire \register_file[11][15] ;
 wire \register_file[11][16] ;
 wire \register_file[11][17] ;
 wire \register_file[11][18] ;
 wire \register_file[11][19] ;
 wire \register_file[11][1] ;
 wire \register_file[11][20] ;
 wire \register_file[11][21] ;
 wire \register_file[11][22] ;
 wire \register_file[11][23] ;
 wire \register_file[11][24] ;
 wire \register_file[11][25] ;
 wire \register_file[11][26] ;
 wire \register_file[11][27] ;
 wire \register_file[11][28] ;
 wire \register_file[11][29] ;
 wire \register_file[11][2] ;
 wire \register_file[11][30] ;
 wire \register_file[11][31] ;
 wire \register_file[11][3] ;
 wire \register_file[11][4] ;
 wire \register_file[11][5] ;
 wire \register_file[11][6] ;
 wire \register_file[11][7] ;
 wire \register_file[11][8] ;
 wire \register_file[11][9] ;
 wire \register_file[12][0] ;
 wire \register_file[12][10] ;
 wire \register_file[12][11] ;
 wire \register_file[12][12] ;
 wire \register_file[12][13] ;
 wire \register_file[12][14] ;
 wire \register_file[12][15] ;
 wire \register_file[12][16] ;
 wire \register_file[12][17] ;
 wire \register_file[12][18] ;
 wire \register_file[12][19] ;
 wire \register_file[12][1] ;
 wire \register_file[12][20] ;
 wire \register_file[12][21] ;
 wire \register_file[12][22] ;
 wire \register_file[12][23] ;
 wire \register_file[12][24] ;
 wire \register_file[12][25] ;
 wire \register_file[12][26] ;
 wire \register_file[12][27] ;
 wire \register_file[12][28] ;
 wire \register_file[12][29] ;
 wire \register_file[12][2] ;
 wire \register_file[12][30] ;
 wire \register_file[12][31] ;
 wire \register_file[12][3] ;
 wire \register_file[12][4] ;
 wire \register_file[12][5] ;
 wire \register_file[12][6] ;
 wire \register_file[12][7] ;
 wire \register_file[12][8] ;
 wire \register_file[12][9] ;
 wire \register_file[13][0] ;
 wire \register_file[13][10] ;
 wire \register_file[13][11] ;
 wire \register_file[13][12] ;
 wire \register_file[13][13] ;
 wire \register_file[13][14] ;
 wire \register_file[13][15] ;
 wire \register_file[13][16] ;
 wire \register_file[13][17] ;
 wire \register_file[13][18] ;
 wire \register_file[13][19] ;
 wire \register_file[13][1] ;
 wire \register_file[13][20] ;
 wire \register_file[13][21] ;
 wire \register_file[13][22] ;
 wire \register_file[13][23] ;
 wire \register_file[13][24] ;
 wire \register_file[13][25] ;
 wire \register_file[13][26] ;
 wire \register_file[13][27] ;
 wire \register_file[13][28] ;
 wire \register_file[13][29] ;
 wire \register_file[13][2] ;
 wire \register_file[13][30] ;
 wire \register_file[13][31] ;
 wire \register_file[13][3] ;
 wire \register_file[13][4] ;
 wire \register_file[13][5] ;
 wire \register_file[13][6] ;
 wire \register_file[13][7] ;
 wire \register_file[13][8] ;
 wire \register_file[13][9] ;
 wire \register_file[14][0] ;
 wire \register_file[14][10] ;
 wire \register_file[14][11] ;
 wire \register_file[14][12] ;
 wire \register_file[14][13] ;
 wire \register_file[14][14] ;
 wire \register_file[14][15] ;
 wire \register_file[14][16] ;
 wire \register_file[14][17] ;
 wire \register_file[14][18] ;
 wire \register_file[14][19] ;
 wire \register_file[14][1] ;
 wire \register_file[14][20] ;
 wire \register_file[14][21] ;
 wire \register_file[14][22] ;
 wire \register_file[14][23] ;
 wire \register_file[14][24] ;
 wire \register_file[14][25] ;
 wire \register_file[14][26] ;
 wire \register_file[14][27] ;
 wire \register_file[14][28] ;
 wire \register_file[14][29] ;
 wire \register_file[14][2] ;
 wire \register_file[14][30] ;
 wire \register_file[14][31] ;
 wire \register_file[14][3] ;
 wire \register_file[14][4] ;
 wire \register_file[14][5] ;
 wire \register_file[14][6] ;
 wire \register_file[14][7] ;
 wire \register_file[14][8] ;
 wire \register_file[14][9] ;
 wire \register_file[15][0] ;
 wire \register_file[15][10] ;
 wire \register_file[15][11] ;
 wire \register_file[15][12] ;
 wire \register_file[15][13] ;
 wire \register_file[15][14] ;
 wire \register_file[15][15] ;
 wire \register_file[15][16] ;
 wire \register_file[15][17] ;
 wire \register_file[15][18] ;
 wire \register_file[15][19] ;
 wire \register_file[15][1] ;
 wire \register_file[15][20] ;
 wire \register_file[15][21] ;
 wire \register_file[15][22] ;
 wire \register_file[15][23] ;
 wire \register_file[15][24] ;
 wire \register_file[15][25] ;
 wire \register_file[15][26] ;
 wire \register_file[15][27] ;
 wire \register_file[15][28] ;
 wire \register_file[15][29] ;
 wire \register_file[15][2] ;
 wire \register_file[15][30] ;
 wire \register_file[15][31] ;
 wire \register_file[15][3] ;
 wire \register_file[15][4] ;
 wire \register_file[15][5] ;
 wire \register_file[15][6] ;
 wire \register_file[15][7] ;
 wire \register_file[15][8] ;
 wire \register_file[15][9] ;
 wire \register_file[16][0] ;
 wire \register_file[16][10] ;
 wire \register_file[16][11] ;
 wire \register_file[16][12] ;
 wire \register_file[16][13] ;
 wire \register_file[16][14] ;
 wire \register_file[16][15] ;
 wire \register_file[16][16] ;
 wire \register_file[16][17] ;
 wire \register_file[16][18] ;
 wire \register_file[16][19] ;
 wire \register_file[16][1] ;
 wire \register_file[16][20] ;
 wire \register_file[16][21] ;
 wire \register_file[16][22] ;
 wire \register_file[16][23] ;
 wire \register_file[16][24] ;
 wire \register_file[16][25] ;
 wire \register_file[16][26] ;
 wire \register_file[16][27] ;
 wire \register_file[16][28] ;
 wire \register_file[16][29] ;
 wire \register_file[16][2] ;
 wire \register_file[16][30] ;
 wire \register_file[16][31] ;
 wire \register_file[16][3] ;
 wire \register_file[16][4] ;
 wire \register_file[16][5] ;
 wire \register_file[16][6] ;
 wire \register_file[16][7] ;
 wire \register_file[16][8] ;
 wire \register_file[16][9] ;
 wire \register_file[17][0] ;
 wire \register_file[17][10] ;
 wire \register_file[17][11] ;
 wire \register_file[17][12] ;
 wire \register_file[17][13] ;
 wire \register_file[17][14] ;
 wire \register_file[17][15] ;
 wire \register_file[17][16] ;
 wire \register_file[17][17] ;
 wire \register_file[17][18] ;
 wire \register_file[17][19] ;
 wire \register_file[17][1] ;
 wire \register_file[17][20] ;
 wire \register_file[17][21] ;
 wire \register_file[17][22] ;
 wire \register_file[17][23] ;
 wire \register_file[17][24] ;
 wire \register_file[17][25] ;
 wire \register_file[17][26] ;
 wire \register_file[17][27] ;
 wire \register_file[17][28] ;
 wire \register_file[17][29] ;
 wire \register_file[17][2] ;
 wire \register_file[17][30] ;
 wire \register_file[17][31] ;
 wire \register_file[17][3] ;
 wire \register_file[17][4] ;
 wire \register_file[17][5] ;
 wire \register_file[17][6] ;
 wire \register_file[17][7] ;
 wire \register_file[17][8] ;
 wire \register_file[17][9] ;
 wire \register_file[18][0] ;
 wire \register_file[18][10] ;
 wire \register_file[18][11] ;
 wire \register_file[18][12] ;
 wire \register_file[18][13] ;
 wire \register_file[18][14] ;
 wire \register_file[18][15] ;
 wire \register_file[18][16] ;
 wire \register_file[18][17] ;
 wire \register_file[18][18] ;
 wire \register_file[18][19] ;
 wire \register_file[18][1] ;
 wire \register_file[18][20] ;
 wire \register_file[18][21] ;
 wire \register_file[18][22] ;
 wire \register_file[18][23] ;
 wire \register_file[18][24] ;
 wire \register_file[18][25] ;
 wire \register_file[18][26] ;
 wire \register_file[18][27] ;
 wire \register_file[18][28] ;
 wire \register_file[18][29] ;
 wire \register_file[18][2] ;
 wire \register_file[18][30] ;
 wire \register_file[18][31] ;
 wire \register_file[18][3] ;
 wire \register_file[18][4] ;
 wire \register_file[18][5] ;
 wire \register_file[18][6] ;
 wire \register_file[18][7] ;
 wire \register_file[18][8] ;
 wire \register_file[18][9] ;
 wire \register_file[19][0] ;
 wire \register_file[19][10] ;
 wire \register_file[19][11] ;
 wire \register_file[19][12] ;
 wire \register_file[19][13] ;
 wire \register_file[19][14] ;
 wire \register_file[19][15] ;
 wire \register_file[19][16] ;
 wire \register_file[19][17] ;
 wire \register_file[19][18] ;
 wire \register_file[19][19] ;
 wire \register_file[19][1] ;
 wire \register_file[19][20] ;
 wire \register_file[19][21] ;
 wire \register_file[19][22] ;
 wire \register_file[19][23] ;
 wire \register_file[19][24] ;
 wire \register_file[19][25] ;
 wire \register_file[19][26] ;
 wire \register_file[19][27] ;
 wire \register_file[19][28] ;
 wire \register_file[19][29] ;
 wire \register_file[19][2] ;
 wire \register_file[19][30] ;
 wire \register_file[19][31] ;
 wire \register_file[19][3] ;
 wire \register_file[19][4] ;
 wire \register_file[19][5] ;
 wire \register_file[19][6] ;
 wire \register_file[19][7] ;
 wire \register_file[19][8] ;
 wire \register_file[19][9] ;
 wire \register_file[1][0] ;
 wire \register_file[1][10] ;
 wire \register_file[1][11] ;
 wire \register_file[1][12] ;
 wire \register_file[1][13] ;
 wire \register_file[1][14] ;
 wire \register_file[1][15] ;
 wire \register_file[1][16] ;
 wire \register_file[1][17] ;
 wire \register_file[1][18] ;
 wire \register_file[1][19] ;
 wire \register_file[1][1] ;
 wire \register_file[1][20] ;
 wire \register_file[1][21] ;
 wire \register_file[1][22] ;
 wire \register_file[1][23] ;
 wire \register_file[1][24] ;
 wire \register_file[1][25] ;
 wire \register_file[1][26] ;
 wire \register_file[1][27] ;
 wire \register_file[1][28] ;
 wire \register_file[1][29] ;
 wire \register_file[1][2] ;
 wire \register_file[1][30] ;
 wire \register_file[1][31] ;
 wire \register_file[1][3] ;
 wire \register_file[1][4] ;
 wire \register_file[1][5] ;
 wire \register_file[1][6] ;
 wire \register_file[1][7] ;
 wire \register_file[1][8] ;
 wire \register_file[1][9] ;
 wire \register_file[20][0] ;
 wire \register_file[20][10] ;
 wire \register_file[20][11] ;
 wire \register_file[20][12] ;
 wire \register_file[20][13] ;
 wire \register_file[20][14] ;
 wire \register_file[20][15] ;
 wire \register_file[20][16] ;
 wire \register_file[20][17] ;
 wire \register_file[20][18] ;
 wire \register_file[20][19] ;
 wire \register_file[20][1] ;
 wire \register_file[20][20] ;
 wire \register_file[20][21] ;
 wire \register_file[20][22] ;
 wire \register_file[20][23] ;
 wire \register_file[20][24] ;
 wire \register_file[20][25] ;
 wire \register_file[20][26] ;
 wire \register_file[20][27] ;
 wire \register_file[20][28] ;
 wire \register_file[20][29] ;
 wire \register_file[20][2] ;
 wire \register_file[20][30] ;
 wire \register_file[20][31] ;
 wire \register_file[20][3] ;
 wire \register_file[20][4] ;
 wire \register_file[20][5] ;
 wire \register_file[20][6] ;
 wire \register_file[20][7] ;
 wire \register_file[20][8] ;
 wire \register_file[20][9] ;
 wire \register_file[21][0] ;
 wire \register_file[21][10] ;
 wire \register_file[21][11] ;
 wire \register_file[21][12] ;
 wire \register_file[21][13] ;
 wire \register_file[21][14] ;
 wire \register_file[21][15] ;
 wire \register_file[21][16] ;
 wire \register_file[21][17] ;
 wire \register_file[21][18] ;
 wire \register_file[21][19] ;
 wire \register_file[21][1] ;
 wire \register_file[21][20] ;
 wire \register_file[21][21] ;
 wire \register_file[21][22] ;
 wire \register_file[21][23] ;
 wire \register_file[21][24] ;
 wire \register_file[21][25] ;
 wire \register_file[21][26] ;
 wire \register_file[21][27] ;
 wire \register_file[21][28] ;
 wire \register_file[21][29] ;
 wire \register_file[21][2] ;
 wire \register_file[21][30] ;
 wire \register_file[21][31] ;
 wire \register_file[21][3] ;
 wire \register_file[21][4] ;
 wire \register_file[21][5] ;
 wire \register_file[21][6] ;
 wire \register_file[21][7] ;
 wire \register_file[21][8] ;
 wire \register_file[21][9] ;
 wire \register_file[22][0] ;
 wire \register_file[22][10] ;
 wire \register_file[22][11] ;
 wire \register_file[22][12] ;
 wire \register_file[22][13] ;
 wire \register_file[22][14] ;
 wire \register_file[22][15] ;
 wire \register_file[22][16] ;
 wire \register_file[22][17] ;
 wire \register_file[22][18] ;
 wire \register_file[22][19] ;
 wire \register_file[22][1] ;
 wire \register_file[22][20] ;
 wire \register_file[22][21] ;
 wire \register_file[22][22] ;
 wire \register_file[22][23] ;
 wire \register_file[22][24] ;
 wire \register_file[22][25] ;
 wire \register_file[22][26] ;
 wire \register_file[22][27] ;
 wire \register_file[22][28] ;
 wire \register_file[22][29] ;
 wire \register_file[22][2] ;
 wire \register_file[22][30] ;
 wire \register_file[22][31] ;
 wire \register_file[22][3] ;
 wire \register_file[22][4] ;
 wire \register_file[22][5] ;
 wire \register_file[22][6] ;
 wire \register_file[22][7] ;
 wire \register_file[22][8] ;
 wire \register_file[22][9] ;
 wire \register_file[23][0] ;
 wire \register_file[23][10] ;
 wire \register_file[23][11] ;
 wire \register_file[23][12] ;
 wire \register_file[23][13] ;
 wire \register_file[23][14] ;
 wire \register_file[23][15] ;
 wire \register_file[23][16] ;
 wire \register_file[23][17] ;
 wire \register_file[23][18] ;
 wire \register_file[23][19] ;
 wire \register_file[23][1] ;
 wire \register_file[23][20] ;
 wire \register_file[23][21] ;
 wire \register_file[23][22] ;
 wire \register_file[23][23] ;
 wire \register_file[23][24] ;
 wire \register_file[23][25] ;
 wire \register_file[23][26] ;
 wire \register_file[23][27] ;
 wire \register_file[23][28] ;
 wire \register_file[23][29] ;
 wire \register_file[23][2] ;
 wire \register_file[23][30] ;
 wire \register_file[23][31] ;
 wire \register_file[23][3] ;
 wire \register_file[23][4] ;
 wire \register_file[23][5] ;
 wire \register_file[23][6] ;
 wire \register_file[23][7] ;
 wire \register_file[23][8] ;
 wire \register_file[23][9] ;
 wire \register_file[24][0] ;
 wire \register_file[24][10] ;
 wire \register_file[24][11] ;
 wire \register_file[24][12] ;
 wire \register_file[24][13] ;
 wire \register_file[24][14] ;
 wire \register_file[24][15] ;
 wire \register_file[24][16] ;
 wire \register_file[24][17] ;
 wire \register_file[24][18] ;
 wire \register_file[24][19] ;
 wire \register_file[24][1] ;
 wire \register_file[24][20] ;
 wire \register_file[24][21] ;
 wire \register_file[24][22] ;
 wire \register_file[24][23] ;
 wire \register_file[24][24] ;
 wire \register_file[24][25] ;
 wire \register_file[24][26] ;
 wire \register_file[24][27] ;
 wire \register_file[24][28] ;
 wire \register_file[24][29] ;
 wire \register_file[24][2] ;
 wire \register_file[24][30] ;
 wire \register_file[24][31] ;
 wire \register_file[24][3] ;
 wire \register_file[24][4] ;
 wire \register_file[24][5] ;
 wire \register_file[24][6] ;
 wire \register_file[24][7] ;
 wire \register_file[24][8] ;
 wire \register_file[24][9] ;
 wire \register_file[25][0] ;
 wire \register_file[25][10] ;
 wire \register_file[25][11] ;
 wire \register_file[25][12] ;
 wire \register_file[25][13] ;
 wire \register_file[25][14] ;
 wire \register_file[25][15] ;
 wire \register_file[25][16] ;
 wire \register_file[25][17] ;
 wire \register_file[25][18] ;
 wire \register_file[25][19] ;
 wire \register_file[25][1] ;
 wire \register_file[25][20] ;
 wire \register_file[25][21] ;
 wire \register_file[25][22] ;
 wire \register_file[25][23] ;
 wire \register_file[25][24] ;
 wire \register_file[25][25] ;
 wire \register_file[25][26] ;
 wire \register_file[25][27] ;
 wire \register_file[25][28] ;
 wire \register_file[25][29] ;
 wire \register_file[25][2] ;
 wire \register_file[25][30] ;
 wire \register_file[25][31] ;
 wire \register_file[25][3] ;
 wire \register_file[25][4] ;
 wire \register_file[25][5] ;
 wire \register_file[25][6] ;
 wire \register_file[25][7] ;
 wire \register_file[25][8] ;
 wire \register_file[25][9] ;
 wire \register_file[26][0] ;
 wire \register_file[26][10] ;
 wire \register_file[26][11] ;
 wire \register_file[26][12] ;
 wire \register_file[26][13] ;
 wire \register_file[26][14] ;
 wire \register_file[26][15] ;
 wire \register_file[26][16] ;
 wire \register_file[26][17] ;
 wire \register_file[26][18] ;
 wire \register_file[26][19] ;
 wire \register_file[26][1] ;
 wire \register_file[26][20] ;
 wire \register_file[26][21] ;
 wire \register_file[26][22] ;
 wire \register_file[26][23] ;
 wire \register_file[26][24] ;
 wire \register_file[26][25] ;
 wire \register_file[26][26] ;
 wire \register_file[26][27] ;
 wire \register_file[26][28] ;
 wire \register_file[26][29] ;
 wire \register_file[26][2] ;
 wire \register_file[26][30] ;
 wire \register_file[26][31] ;
 wire \register_file[26][3] ;
 wire \register_file[26][4] ;
 wire \register_file[26][5] ;
 wire \register_file[26][6] ;
 wire \register_file[26][7] ;
 wire \register_file[26][8] ;
 wire \register_file[26][9] ;
 wire \register_file[27][0] ;
 wire \register_file[27][10] ;
 wire \register_file[27][11] ;
 wire \register_file[27][12] ;
 wire \register_file[27][13] ;
 wire \register_file[27][14] ;
 wire \register_file[27][15] ;
 wire \register_file[27][16] ;
 wire \register_file[27][17] ;
 wire \register_file[27][18] ;
 wire \register_file[27][19] ;
 wire \register_file[27][1] ;
 wire \register_file[27][20] ;
 wire \register_file[27][21] ;
 wire \register_file[27][22] ;
 wire \register_file[27][23] ;
 wire \register_file[27][24] ;
 wire \register_file[27][25] ;
 wire \register_file[27][26] ;
 wire \register_file[27][27] ;
 wire \register_file[27][28] ;
 wire \register_file[27][29] ;
 wire \register_file[27][2] ;
 wire \register_file[27][30] ;
 wire \register_file[27][31] ;
 wire \register_file[27][3] ;
 wire \register_file[27][4] ;
 wire \register_file[27][5] ;
 wire \register_file[27][6] ;
 wire \register_file[27][7] ;
 wire \register_file[27][8] ;
 wire \register_file[27][9] ;
 wire \register_file[28][0] ;
 wire \register_file[28][10] ;
 wire \register_file[28][11] ;
 wire \register_file[28][12] ;
 wire \register_file[28][13] ;
 wire \register_file[28][14] ;
 wire \register_file[28][15] ;
 wire \register_file[28][16] ;
 wire \register_file[28][17] ;
 wire \register_file[28][18] ;
 wire \register_file[28][19] ;
 wire \register_file[28][1] ;
 wire \register_file[28][20] ;
 wire \register_file[28][21] ;
 wire \register_file[28][22] ;
 wire \register_file[28][23] ;
 wire \register_file[28][24] ;
 wire \register_file[28][25] ;
 wire \register_file[28][26] ;
 wire \register_file[28][27] ;
 wire \register_file[28][28] ;
 wire \register_file[28][29] ;
 wire \register_file[28][2] ;
 wire \register_file[28][30] ;
 wire \register_file[28][31] ;
 wire \register_file[28][3] ;
 wire \register_file[28][4] ;
 wire \register_file[28][5] ;
 wire \register_file[28][6] ;
 wire \register_file[28][7] ;
 wire \register_file[28][8] ;
 wire \register_file[28][9] ;
 wire \register_file[29][0] ;
 wire \register_file[29][10] ;
 wire \register_file[29][11] ;
 wire \register_file[29][12] ;
 wire \register_file[29][13] ;
 wire \register_file[29][14] ;
 wire \register_file[29][15] ;
 wire \register_file[29][16] ;
 wire \register_file[29][17] ;
 wire \register_file[29][18] ;
 wire \register_file[29][19] ;
 wire \register_file[29][1] ;
 wire \register_file[29][20] ;
 wire \register_file[29][21] ;
 wire \register_file[29][22] ;
 wire \register_file[29][23] ;
 wire \register_file[29][24] ;
 wire \register_file[29][25] ;
 wire \register_file[29][26] ;
 wire \register_file[29][27] ;
 wire \register_file[29][28] ;
 wire \register_file[29][29] ;
 wire \register_file[29][2] ;
 wire \register_file[29][30] ;
 wire \register_file[29][31] ;
 wire \register_file[29][3] ;
 wire \register_file[29][4] ;
 wire \register_file[29][5] ;
 wire \register_file[29][6] ;
 wire \register_file[29][7] ;
 wire \register_file[29][8] ;
 wire \register_file[29][9] ;
 wire \register_file[2][0] ;
 wire \register_file[2][10] ;
 wire \register_file[2][11] ;
 wire \register_file[2][12] ;
 wire \register_file[2][13] ;
 wire \register_file[2][14] ;
 wire \register_file[2][15] ;
 wire \register_file[2][16] ;
 wire \register_file[2][17] ;
 wire \register_file[2][18] ;
 wire \register_file[2][19] ;
 wire \register_file[2][1] ;
 wire \register_file[2][20] ;
 wire \register_file[2][21] ;
 wire \register_file[2][22] ;
 wire \register_file[2][23] ;
 wire \register_file[2][24] ;
 wire \register_file[2][25] ;
 wire \register_file[2][26] ;
 wire \register_file[2][27] ;
 wire \register_file[2][28] ;
 wire \register_file[2][29] ;
 wire \register_file[2][2] ;
 wire \register_file[2][30] ;
 wire \register_file[2][31] ;
 wire \register_file[2][3] ;
 wire \register_file[2][4] ;
 wire \register_file[2][5] ;
 wire \register_file[2][6] ;
 wire \register_file[2][7] ;
 wire \register_file[2][8] ;
 wire \register_file[2][9] ;
 wire \register_file[30][0] ;
 wire \register_file[30][10] ;
 wire \register_file[30][11] ;
 wire \register_file[30][12] ;
 wire \register_file[30][13] ;
 wire \register_file[30][14] ;
 wire \register_file[30][15] ;
 wire \register_file[30][16] ;
 wire \register_file[30][17] ;
 wire \register_file[30][18] ;
 wire \register_file[30][19] ;
 wire \register_file[30][1] ;
 wire \register_file[30][20] ;
 wire \register_file[30][21] ;
 wire \register_file[30][22] ;
 wire \register_file[30][23] ;
 wire \register_file[30][24] ;
 wire \register_file[30][25] ;
 wire \register_file[30][26] ;
 wire \register_file[30][27] ;
 wire \register_file[30][28] ;
 wire \register_file[30][29] ;
 wire \register_file[30][2] ;
 wire \register_file[30][30] ;
 wire \register_file[30][31] ;
 wire \register_file[30][3] ;
 wire \register_file[30][4] ;
 wire \register_file[30][5] ;
 wire \register_file[30][6] ;
 wire \register_file[30][7] ;
 wire \register_file[30][8] ;
 wire \register_file[30][9] ;
 wire \register_file[31][0] ;
 wire \register_file[31][10] ;
 wire \register_file[31][11] ;
 wire \register_file[31][12] ;
 wire \register_file[31][13] ;
 wire \register_file[31][14] ;
 wire \register_file[31][15] ;
 wire \register_file[31][16] ;
 wire \register_file[31][17] ;
 wire \register_file[31][18] ;
 wire \register_file[31][19] ;
 wire \register_file[31][1] ;
 wire \register_file[31][20] ;
 wire \register_file[31][21] ;
 wire \register_file[31][22] ;
 wire \register_file[31][23] ;
 wire \register_file[31][24] ;
 wire \register_file[31][25] ;
 wire \register_file[31][26] ;
 wire \register_file[31][27] ;
 wire \register_file[31][28] ;
 wire \register_file[31][29] ;
 wire \register_file[31][2] ;
 wire \register_file[31][30] ;
 wire \register_file[31][31] ;
 wire \register_file[31][3] ;
 wire \register_file[31][4] ;
 wire \register_file[31][5] ;
 wire \register_file[31][6] ;
 wire \register_file[31][7] ;
 wire \register_file[31][8] ;
 wire \register_file[31][9] ;
 wire \register_file[3][0] ;
 wire \register_file[3][10] ;
 wire \register_file[3][11] ;
 wire \register_file[3][12] ;
 wire \register_file[3][13] ;
 wire \register_file[3][14] ;
 wire \register_file[3][15] ;
 wire \register_file[3][16] ;
 wire \register_file[3][17] ;
 wire \register_file[3][18] ;
 wire \register_file[3][19] ;
 wire \register_file[3][1] ;
 wire \register_file[3][20] ;
 wire \register_file[3][21] ;
 wire \register_file[3][22] ;
 wire \register_file[3][23] ;
 wire \register_file[3][24] ;
 wire \register_file[3][25] ;
 wire \register_file[3][26] ;
 wire \register_file[3][27] ;
 wire \register_file[3][28] ;
 wire \register_file[3][29] ;
 wire \register_file[3][2] ;
 wire \register_file[3][30] ;
 wire \register_file[3][31] ;
 wire \register_file[3][3] ;
 wire \register_file[3][4] ;
 wire \register_file[3][5] ;
 wire \register_file[3][6] ;
 wire \register_file[3][7] ;
 wire \register_file[3][8] ;
 wire \register_file[3][9] ;
 wire \register_file[4][0] ;
 wire \register_file[4][10] ;
 wire \register_file[4][11] ;
 wire \register_file[4][12] ;
 wire \register_file[4][13] ;
 wire \register_file[4][14] ;
 wire \register_file[4][15] ;
 wire \register_file[4][16] ;
 wire \register_file[4][17] ;
 wire \register_file[4][18] ;
 wire \register_file[4][19] ;
 wire \register_file[4][1] ;
 wire \register_file[4][20] ;
 wire \register_file[4][21] ;
 wire \register_file[4][22] ;
 wire \register_file[4][23] ;
 wire \register_file[4][24] ;
 wire \register_file[4][25] ;
 wire \register_file[4][26] ;
 wire \register_file[4][27] ;
 wire \register_file[4][28] ;
 wire \register_file[4][29] ;
 wire \register_file[4][2] ;
 wire \register_file[4][30] ;
 wire \register_file[4][31] ;
 wire \register_file[4][3] ;
 wire \register_file[4][4] ;
 wire \register_file[4][5] ;
 wire \register_file[4][6] ;
 wire \register_file[4][7] ;
 wire \register_file[4][8] ;
 wire \register_file[4][9] ;
 wire \register_file[5][0] ;
 wire \register_file[5][10] ;
 wire \register_file[5][11] ;
 wire \register_file[5][12] ;
 wire \register_file[5][13] ;
 wire \register_file[5][14] ;
 wire \register_file[5][15] ;
 wire \register_file[5][16] ;
 wire \register_file[5][17] ;
 wire \register_file[5][18] ;
 wire \register_file[5][19] ;
 wire \register_file[5][1] ;
 wire \register_file[5][20] ;
 wire \register_file[5][21] ;
 wire \register_file[5][22] ;
 wire \register_file[5][23] ;
 wire \register_file[5][24] ;
 wire \register_file[5][25] ;
 wire \register_file[5][26] ;
 wire \register_file[5][27] ;
 wire \register_file[5][28] ;
 wire \register_file[5][29] ;
 wire \register_file[5][2] ;
 wire \register_file[5][30] ;
 wire \register_file[5][31] ;
 wire \register_file[5][3] ;
 wire \register_file[5][4] ;
 wire \register_file[5][5] ;
 wire \register_file[5][6] ;
 wire \register_file[5][7] ;
 wire \register_file[5][8] ;
 wire \register_file[5][9] ;
 wire \register_file[6][0] ;
 wire \register_file[6][10] ;
 wire \register_file[6][11] ;
 wire \register_file[6][12] ;
 wire \register_file[6][13] ;
 wire \register_file[6][14] ;
 wire \register_file[6][15] ;
 wire \register_file[6][16] ;
 wire \register_file[6][17] ;
 wire \register_file[6][18] ;
 wire \register_file[6][19] ;
 wire \register_file[6][1] ;
 wire \register_file[6][20] ;
 wire \register_file[6][21] ;
 wire \register_file[6][22] ;
 wire \register_file[6][23] ;
 wire \register_file[6][24] ;
 wire \register_file[6][25] ;
 wire \register_file[6][26] ;
 wire \register_file[6][27] ;
 wire \register_file[6][28] ;
 wire \register_file[6][29] ;
 wire \register_file[6][2] ;
 wire \register_file[6][30] ;
 wire \register_file[6][31] ;
 wire \register_file[6][3] ;
 wire \register_file[6][4] ;
 wire \register_file[6][5] ;
 wire \register_file[6][6] ;
 wire \register_file[6][7] ;
 wire \register_file[6][8] ;
 wire \register_file[6][9] ;
 wire \register_file[7][0] ;
 wire \register_file[7][10] ;
 wire \register_file[7][11] ;
 wire \register_file[7][12] ;
 wire \register_file[7][13] ;
 wire \register_file[7][14] ;
 wire \register_file[7][15] ;
 wire \register_file[7][16] ;
 wire \register_file[7][17] ;
 wire \register_file[7][18] ;
 wire \register_file[7][19] ;
 wire \register_file[7][1] ;
 wire \register_file[7][20] ;
 wire \register_file[7][21] ;
 wire \register_file[7][22] ;
 wire \register_file[7][23] ;
 wire \register_file[7][24] ;
 wire \register_file[7][25] ;
 wire \register_file[7][26] ;
 wire \register_file[7][27] ;
 wire \register_file[7][28] ;
 wire \register_file[7][29] ;
 wire \register_file[7][2] ;
 wire \register_file[7][30] ;
 wire \register_file[7][31] ;
 wire \register_file[7][3] ;
 wire \register_file[7][4] ;
 wire \register_file[7][5] ;
 wire \register_file[7][6] ;
 wire \register_file[7][7] ;
 wire \register_file[7][8] ;
 wire \register_file[7][9] ;
 wire \register_file[8][0] ;
 wire \register_file[8][10] ;
 wire \register_file[8][11] ;
 wire \register_file[8][12] ;
 wire \register_file[8][13] ;
 wire \register_file[8][14] ;
 wire \register_file[8][15] ;
 wire \register_file[8][16] ;
 wire \register_file[8][17] ;
 wire \register_file[8][18] ;
 wire \register_file[8][19] ;
 wire \register_file[8][1] ;
 wire \register_file[8][20] ;
 wire \register_file[8][21] ;
 wire \register_file[8][22] ;
 wire \register_file[8][23] ;
 wire \register_file[8][24] ;
 wire \register_file[8][25] ;
 wire \register_file[8][26] ;
 wire \register_file[8][27] ;
 wire \register_file[8][28] ;
 wire \register_file[8][29] ;
 wire \register_file[8][2] ;
 wire \register_file[8][30] ;
 wire \register_file[8][31] ;
 wire \register_file[8][3] ;
 wire \register_file[8][4] ;
 wire \register_file[8][5] ;
 wire \register_file[8][6] ;
 wire \register_file[8][7] ;
 wire \register_file[8][8] ;
 wire \register_file[8][9] ;
 wire \register_file[9][0] ;
 wire \register_file[9][10] ;
 wire \register_file[9][11] ;
 wire \register_file[9][12] ;
 wire \register_file[9][13] ;
 wire \register_file[9][14] ;
 wire \register_file[9][15] ;
 wire \register_file[9][16] ;
 wire \register_file[9][17] ;
 wire \register_file[9][18] ;
 wire \register_file[9][19] ;
 wire \register_file[9][1] ;
 wire \register_file[9][20] ;
 wire \register_file[9][21] ;
 wire \register_file[9][22] ;
 wire \register_file[9][23] ;
 wire \register_file[9][24] ;
 wire \register_file[9][25] ;
 wire \register_file[9][26] ;
 wire \register_file[9][27] ;
 wire \register_file[9][28] ;
 wire \register_file[9][29] ;
 wire \register_file[9][2] ;
 wire \register_file[9][30] ;
 wire \register_file[9][31] ;
 wire \register_file[9][3] ;
 wire \register_file[9][4] ;
 wire \register_file[9][5] ;
 wire \register_file[9][6] ;
 wire \register_file[9][7] ;
 wire \register_file[9][8] ;
 wire \register_file[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07774_ (.A1(_03105_),
    .A2(_03109_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07775_ (.A1(_02940_),
    .A2(\register_file[12][23] ),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07776_ (.A1(_03027_),
    .A2(\register_file[13][23] ),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07777_ (.A1(_03111_),
    .A2(_03026_),
    .A3(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07778_ (.A1(_02857_),
    .A2(\register_file[14][23] ),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07779_ (.A1(_02859_),
    .A2(\register_file[15][23] ),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07780_ (.A1(_03114_),
    .A2(_02945_),
    .A3(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07781_ (.A1(_03113_),
    .A2(_03116_),
    .A3(_02862_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07782_ (.A1(_03110_),
    .A2(_03117_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07783_ (.A1(_02865_),
    .A2(\register_file[6][23] ),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07784_ (.I(\register_file[7][23] ),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07785_ (.A1(_03120_),
    .A2(_03037_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07786_ (.A1(_03119_),
    .A2(_03121_),
    .A3(_02953_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07787_ (.I(\register_file[4][23] ),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07788_ (.A1(_02786_),
    .A2(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07789_ (.I(\register_file[5][23] ),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07790_ (.A1(_03125_),
    .A2(_02958_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07791_ (.A1(_03124_),
    .A2(_03126_),
    .A3(_02960_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07792_ (.A1(_03122_),
    .A2(_03127_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07793_ (.A1(_03128_),
    .A2(_02793_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07794_ (.A1(_02964_),
    .A2(\register_file[2][23] ),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07795_ (.I(\register_file[3][23] ),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07796_ (.I(_01155_),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07797_ (.A1(_03131_),
    .A2(_03132_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07798_ (.A1(_02877_),
    .A2(_03130_),
    .A3(_03133_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07799_ (.A1(_03051_),
    .A2(\register_file[1][23] ),
    .B(_03052_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07800_ (.A1(_03134_),
    .A2(_03135_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07801_ (.I(_03136_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07802_ (.A1(_03129_),
    .A2(_03137_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07803_ (.A1(_03118_),
    .A2(_03138_),
    .A3(_02886_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07804_ (.A1(_03098_),
    .A2(_03139_),
    .B(_02888_),
    .ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07805_ (.A1(_02889_),
    .A2(\register_file[16][24] ),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07806_ (.A1(_02805_),
    .A2(\register_file[17][24] ),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07807_ (.A1(_03140_),
    .A2(_03141_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07808_ (.A1(_03142_),
    .A2(_02808_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07809_ (.A1(_03143_),
    .A2(_02978_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07810_ (.A1(_03063_),
    .A2(\register_file[19][24] ),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07811_ (.A1(_02812_),
    .A2(\register_file[18][24] ),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07812_ (.A1(_03145_),
    .A2(_03146_),
    .B(_02814_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07813_ (.A1(_03144_),
    .A2(_03147_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07814_ (.A1(_03068_),
    .A2(\register_file[20][24] ),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07815_ (.I(_01083_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07816_ (.A1(_02818_),
    .A2(\register_file[21][24] ),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07817_ (.A1(_03149_),
    .A2(_03150_),
    .A3(_03151_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07818_ (.I(_01071_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07819_ (.A1(_03153_),
    .A2(\register_file[22][24] ),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07820_ (.I(_01325_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07821_ (.A1(_02903_),
    .A2(\register_file[23][24] ),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07822_ (.A1(_03154_),
    .A2(_03155_),
    .A3(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07823_ (.A1(_03152_),
    .A2(_03157_),
    .A3(_03075_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07824_ (.A1(_03148_),
    .A2(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07825_ (.A1(_02826_),
    .A2(\register_file[24][24] ),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07826_ (.A1(_02993_),
    .A2(\register_file[25][24] ),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07827_ (.A1(_03160_),
    .A2(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07828_ (.I(_01114_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07829_ (.A1(_03162_),
    .A2(_03163_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07830_ (.A1(_03164_),
    .A2(_02912_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07831_ (.A1(_02998_),
    .A2(\register_file[27][24] ),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07832_ (.A1(_03084_),
    .A2(\register_file[26][24] ),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07833_ (.I(_01125_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07834_ (.A1(_03166_),
    .A2(_03167_),
    .B(_03168_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07835_ (.A1(_03165_),
    .A2(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07836_ (.A1(_03003_),
    .A2(\register_file[28][24] ),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07837_ (.A1(_03090_),
    .A2(\register_file[29][24] ),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07838_ (.A1(_03171_),
    .A2(_03089_),
    .A3(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07839_ (.A1(_03007_),
    .A2(\register_file[30][24] ),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07840_ (.A1(_03010_),
    .A2(\register_file[31][24] ),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07841_ (.A1(_03174_),
    .A2(_03009_),
    .A3(_03175_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07842_ (.A1(_03173_),
    .A2(_03176_),
    .A3(_02924_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07843_ (.A1(_03170_),
    .A2(_03177_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07844_ (.I(_01104_),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07845_ (.A1(_03159_),
    .A2(_03178_),
    .A3(_03179_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07846_ (.I(_01079_),
    .Z(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07847_ (.A1(_03181_),
    .A2(\register_file[8][24] ),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07848_ (.A1(_02929_),
    .A2(\register_file[9][24] ),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07849_ (.A1(_03182_),
    .A2(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07850_ (.A1(_03184_),
    .A2(_03102_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07851_ (.A1(_03185_),
    .A2(_03104_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07852_ (.A1(_02934_),
    .A2(\register_file[11][24] ),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07853_ (.A1(_02936_),
    .A2(\register_file[10][24] ),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07854_ (.A1(_03187_),
    .A2(_03188_),
    .B(_03108_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07855_ (.A1(_03186_),
    .A2(_03189_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07856_ (.A1(_02940_),
    .A2(\register_file[12][24] ),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07857_ (.A1(_03027_),
    .A2(\register_file[13][24] ),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07858_ (.A1(_03191_),
    .A2(_03026_),
    .A3(_03192_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07859_ (.A1(_02857_),
    .A2(\register_file[14][24] ),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07860_ (.A1(_02859_),
    .A2(\register_file[15][24] ),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07861_ (.A1(_03194_),
    .A2(_02945_),
    .A3(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07862_ (.A1(_03193_),
    .A2(_03196_),
    .A3(_02862_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07863_ (.A1(_03190_),
    .A2(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07864_ (.A1(_02865_),
    .A2(\register_file[6][24] ),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07865_ (.I(\register_file[7][24] ),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07866_ (.A1(_03200_),
    .A2(_03037_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07867_ (.A1(_03199_),
    .A2(_03201_),
    .A3(_02953_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07868_ (.I(_01530_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07869_ (.I(\register_file[4][24] ),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07870_ (.A1(_03203_),
    .A2(_03204_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07871_ (.I(\register_file[5][24] ),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07872_ (.A1(_03206_),
    .A2(_02958_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07873_ (.A1(_03205_),
    .A2(_03207_),
    .A3(_02960_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07874_ (.A1(_03202_),
    .A2(_03208_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07875_ (.I(_01021_),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07876_ (.A1(_03209_),
    .A2(_03210_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07877_ (.A1(_02964_),
    .A2(\register_file[2][24] ),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07878_ (.I(\register_file[3][24] ),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07879_ (.A1(_03213_),
    .A2(_03132_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07880_ (.A1(_02877_),
    .A2(_03212_),
    .A3(_03214_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07881_ (.A1(_03051_),
    .A2(\register_file[1][24] ),
    .B(_03052_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07882_ (.A1(_03215_),
    .A2(_03216_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07883_ (.I(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07884_ (.A1(_03211_),
    .A2(_03218_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07885_ (.A1(_03198_),
    .A2(_03219_),
    .A3(_02886_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07886_ (.A1(_03180_),
    .A2(_03220_),
    .B(_02888_),
    .ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07887_ (.A1(_02889_),
    .A2(\register_file[24][25] ),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07888_ (.I(_01058_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07889_ (.A1(_03222_),
    .A2(\register_file[25][25] ),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07890_ (.A1(_03221_),
    .A2(_03223_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07891_ (.I(_01062_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07892_ (.A1(_03224_),
    .A2(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07893_ (.A1(_03226_),
    .A2(_01066_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07894_ (.A1(_03063_),
    .A2(\register_file[27][25] ),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07895_ (.I(_01042_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07896_ (.A1(_03229_),
    .A2(\register_file[26][25] ),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07897_ (.I(_01559_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07898_ (.A1(_03228_),
    .A2(_03230_),
    .B(_03231_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07899_ (.A1(_03227_),
    .A2(_03232_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07900_ (.A1(_03068_),
    .A2(\register_file[28][25] ),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07901_ (.I(_01085_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07902_ (.A1(_03235_),
    .A2(\register_file[29][25] ),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07903_ (.A1(_03234_),
    .A2(_03150_),
    .A3(_03236_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07904_ (.A1(_03153_),
    .A2(\register_file[30][25] ),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07905_ (.A1(_02903_),
    .A2(\register_file[31][25] ),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07906_ (.A1(_03238_),
    .A2(_03155_),
    .A3(_03239_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07907_ (.A1(_03237_),
    .A2(_03240_),
    .A3(_03075_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07908_ (.A1(_03233_),
    .A2(_03241_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07909_ (.I(_01107_),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07910_ (.A1(_03243_),
    .A2(\register_file[16][25] ),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07911_ (.A1(_02993_),
    .A2(\register_file[17][25] ),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07912_ (.A1(_03244_),
    .A2(_03245_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07913_ (.A1(_03246_),
    .A2(_03163_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07914_ (.A1(_03247_),
    .A2(_01010_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07915_ (.A1(_02998_),
    .A2(\register_file[19][25] ),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07916_ (.A1(_03084_),
    .A2(\register_file[18][25] ),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07917_ (.A1(_03249_),
    .A2(_03250_),
    .B(_03168_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07918_ (.A1(_03248_),
    .A2(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07919_ (.A1(_03003_),
    .A2(\register_file[20][25] ),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07920_ (.A1(_03090_),
    .A2(\register_file[21][25] ),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07921_ (.A1(_03253_),
    .A2(_03089_),
    .A3(_03254_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07922_ (.A1(_03007_),
    .A2(\register_file[22][25] ),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07923_ (.A1(_03010_),
    .A2(\register_file[23][25] ),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07924_ (.A1(_03256_),
    .A2(_03009_),
    .A3(_03257_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07925_ (.A1(_03255_),
    .A2(_03258_),
    .A3(_02924_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07926_ (.A1(_03252_),
    .A2(_03259_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07927_ (.A1(_03242_),
    .A2(_03260_),
    .A3(_03179_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07928_ (.A1(_03181_),
    .A2(\register_file[8][25] ),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07929_ (.A1(_02929_),
    .A2(\register_file[9][25] ),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07930_ (.A1(_03262_),
    .A2(_03263_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07931_ (.A1(_03264_),
    .A2(_03102_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07932_ (.A1(_03265_),
    .A2(_03104_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07933_ (.A1(_02934_),
    .A2(\register_file[11][25] ),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07934_ (.A1(_02936_),
    .A2(\register_file[10][25] ),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07935_ (.A1(_03267_),
    .A2(_03268_),
    .B(_03108_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07936_ (.A1(_03266_),
    .A2(_03269_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07937_ (.A1(_02940_),
    .A2(\register_file[12][25] ),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07938_ (.A1(_03027_),
    .A2(\register_file[13][25] ),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07939_ (.A1(_03271_),
    .A2(_03026_),
    .A3(_03272_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07940_ (.I(_01161_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07941_ (.A1(_03274_),
    .A2(\register_file[14][25] ),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07942_ (.I(_01455_),
    .Z(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07943_ (.A1(_03276_),
    .A2(\register_file[15][25] ),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07944_ (.A1(_03275_),
    .A2(_02945_),
    .A3(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07945_ (.I(_01051_),
    .Z(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07946_ (.A1(_03273_),
    .A2(_03278_),
    .A3(_03279_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07947_ (.A1(_03270_),
    .A2(_03280_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07948_ (.I(_01178_),
    .Z(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07949_ (.A1(_03282_),
    .A2(\register_file[6][25] ),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07950_ (.I(\register_file[7][25] ),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07951_ (.A1(_03284_),
    .A2(_03037_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07952_ (.A1(_03283_),
    .A2(_03285_),
    .A3(_02953_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07953_ (.I(\register_file[4][25] ),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07954_ (.A1(_03203_),
    .A2(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07955_ (.I(\register_file[5][25] ),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07956_ (.A1(_03289_),
    .A2(_02958_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07957_ (.A1(_03288_),
    .A2(_03290_),
    .A3(_02960_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07958_ (.A1(_03286_),
    .A2(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07959_ (.A1(_03292_),
    .A2(_03210_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07960_ (.I(_01175_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07961_ (.A1(_02964_),
    .A2(\register_file[2][25] ),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07962_ (.I(\register_file[3][25] ),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07963_ (.A1(_03296_),
    .A2(_03132_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07964_ (.A1(_03294_),
    .A2(_03295_),
    .A3(_03297_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07965_ (.A1(_03051_),
    .A2(\register_file[1][25] ),
    .B(_03052_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07966_ (.A1(_03298_),
    .A2(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07967_ (.I(_03300_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07968_ (.A1(_03293_),
    .A2(_03301_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07969_ (.I(_01193_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07970_ (.A1(_03281_),
    .A2(_03302_),
    .A3(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07971_ (.I(_01199_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07972_ (.A1(_03261_),
    .A2(_03304_),
    .B(_03305_),
    .ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07973_ (.I(_01055_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07974_ (.A1(_03306_),
    .A2(\register_file[16][26] ),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07975_ (.A1(_03222_),
    .A2(\register_file[17][26] ),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07976_ (.A1(_03307_),
    .A2(_03308_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(_03309_),
    .A2(_03225_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07978_ (.A1(_03310_),
    .A2(_02978_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07979_ (.A1(_03063_),
    .A2(\register_file[19][26] ),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07980_ (.A1(_03229_),
    .A2(\register_file[18][26] ),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07981_ (.A1(_03312_),
    .A2(_03313_),
    .B(_03231_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07982_ (.A1(_03311_),
    .A2(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07983_ (.A1(_03068_),
    .A2(\register_file[20][26] ),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07984_ (.A1(_03235_),
    .A2(\register_file[21][26] ),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07985_ (.A1(_03316_),
    .A2(_03150_),
    .A3(_03317_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07986_ (.A1(_03153_),
    .A2(\register_file[22][26] ),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07987_ (.I(_01649_),
    .Z(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07988_ (.A1(_03320_),
    .A2(\register_file[23][26] ),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07989_ (.A1(_03319_),
    .A2(_03155_),
    .A3(_03321_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07990_ (.A1(_03318_),
    .A2(_03322_),
    .A3(_03075_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07991_ (.A1(_03315_),
    .A2(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07992_ (.A1(_03243_),
    .A2(\register_file[24][26] ),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07993_ (.A1(_02993_),
    .A2(\register_file[25][26] ),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07994_ (.A1(_03325_),
    .A2(_03326_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07995_ (.A1(_03327_),
    .A2(_03163_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07996_ (.A1(_03328_),
    .A2(_02912_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07997_ (.A1(_02998_),
    .A2(\register_file[27][26] ),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07998_ (.A1(_03084_),
    .A2(\register_file[26][26] ),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07999_ (.A1(_03330_),
    .A2(_03331_),
    .B(_03168_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08000_ (.A1(_03329_),
    .A2(_03332_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08001_ (.A1(_03003_),
    .A2(\register_file[28][26] ),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08002_ (.A1(_03090_),
    .A2(\register_file[29][26] ),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08003_ (.A1(_03334_),
    .A2(_03089_),
    .A3(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08004_ (.A1(_03007_),
    .A2(\register_file[30][26] ),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08005_ (.A1(_03010_),
    .A2(\register_file[31][26] ),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08006_ (.A1(_03337_),
    .A2(_03009_),
    .A3(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08007_ (.I(_01670_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08008_ (.A1(_03336_),
    .A2(_03339_),
    .A3(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08009_ (.A1(_03333_),
    .A2(_03341_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08010_ (.A1(_03324_),
    .A2(_03342_),
    .A3(_03179_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08011_ (.A1(_03181_),
    .A2(\register_file[8][26] ),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08012_ (.I(_01013_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08013_ (.A1(_03345_),
    .A2(\register_file[9][26] ),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08014_ (.A1(_03344_),
    .A2(_03346_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08015_ (.A1(_03347_),
    .A2(_03102_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08016_ (.A1(_03348_),
    .A2(_03104_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08017_ (.I(_01681_),
    .Z(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08018_ (.A1(_03350_),
    .A2(\register_file[11][26] ),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08019_ (.I(_01138_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08020_ (.A1(_03352_),
    .A2(\register_file[10][26] ),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08021_ (.A1(_03351_),
    .A2(_03353_),
    .B(_03108_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08022_ (.A1(_03349_),
    .A2(_03354_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08023_ (.I(_01018_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08024_ (.A1(_03356_),
    .A2(\register_file[12][26] ),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08025_ (.A1(_03027_),
    .A2(\register_file[13][26] ),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08026_ (.A1(_03357_),
    .A2(_03026_),
    .A3(_03358_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08027_ (.A1(_03274_),
    .A2(\register_file[14][26] ),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08028_ (.I(_01693_),
    .Z(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08029_ (.A1(_03276_),
    .A2(\register_file[15][26] ),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08030_ (.A1(_03360_),
    .A2(_03361_),
    .A3(_03362_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08031_ (.A1(_03359_),
    .A2(_03363_),
    .A3(_03279_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08032_ (.A1(_03355_),
    .A2(_03364_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08033_ (.A1(_03282_),
    .A2(\register_file[6][26] ),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08034_ (.I(\register_file[7][26] ),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08035_ (.A1(_03367_),
    .A2(_03037_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08036_ (.I(_01092_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08037_ (.A1(_03366_),
    .A2(_03368_),
    .A3(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08038_ (.I(\register_file[4][26] ),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08039_ (.A1(_03203_),
    .A2(_03371_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08040_ (.I(\register_file[5][26] ),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08041_ (.I(_00999_),
    .Z(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08042_ (.A1(_03373_),
    .A2(_03374_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08043_ (.I(_01034_),
    .Z(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08044_ (.A1(_03372_),
    .A2(_03375_),
    .A3(_03376_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08045_ (.A1(_03370_),
    .A2(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08046_ (.A1(_03378_),
    .A2(_03210_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08047_ (.I(_01151_),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08048_ (.A1(_03380_),
    .A2(\register_file[2][26] ),
    .Z(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08049_ (.I(\register_file[3][26] ),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08050_ (.A1(_03382_),
    .A2(_03132_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08051_ (.A1(_03294_),
    .A2(_03381_),
    .A3(_03383_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08052_ (.A1(_03051_),
    .A2(\register_file[1][26] ),
    .B(_03052_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08053_ (.A1(_03384_),
    .A2(_03385_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08054_ (.I(_03386_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08055_ (.A1(_03379_),
    .A2(_03387_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08056_ (.A1(_03365_),
    .A2(_03388_),
    .A3(_03303_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08057_ (.A1(_03343_),
    .A2(_03389_),
    .B(_03305_),
    .ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08058_ (.A1(_03306_),
    .A2(\register_file[16][27] ),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08059_ (.A1(_03222_),
    .A2(\register_file[17][27] ),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08060_ (.A1(_03390_),
    .A2(_03391_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08061_ (.A1(_03392_),
    .A2(_03225_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08062_ (.A1(_03393_),
    .A2(_02978_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(_03063_),
    .A2(\register_file[19][27] ),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08064_ (.A1(_03229_),
    .A2(\register_file[18][27] ),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08065_ (.A1(_03395_),
    .A2(_03396_),
    .B(_03231_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08066_ (.A1(_03394_),
    .A2(_03397_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08067_ (.A1(_03068_),
    .A2(\register_file[20][27] ),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08068_ (.A1(_03235_),
    .A2(\register_file[21][27] ),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08069_ (.A1(_03399_),
    .A2(_03150_),
    .A3(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08070_ (.A1(_03153_),
    .A2(\register_file[22][27] ),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08071_ (.A1(_03320_),
    .A2(\register_file[23][27] ),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08072_ (.A1(_03402_),
    .A2(_03155_),
    .A3(_03403_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08073_ (.A1(_03401_),
    .A2(_03404_),
    .A3(_03075_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08074_ (.A1(_03398_),
    .A2(_03405_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08075_ (.A1(_03243_),
    .A2(\register_file[24][27] ),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08076_ (.A1(_01111_),
    .A2(\register_file[25][27] ),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08077_ (.A1(_03407_),
    .A2(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08078_ (.A1(_03409_),
    .A2(_03163_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08079_ (.A1(_03410_),
    .A2(_02912_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08080_ (.A1(_01120_),
    .A2(\register_file[27][27] ),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08081_ (.A1(_03084_),
    .A2(\register_file[26][27] ),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08082_ (.A1(_03412_),
    .A2(_03413_),
    .B(_03168_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08083_ (.A1(_03411_),
    .A2(_03414_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08084_ (.A1(_01130_),
    .A2(\register_file[28][27] ),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08085_ (.A1(_03090_),
    .A2(\register_file[29][27] ),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08086_ (.A1(_03416_),
    .A2(_03089_),
    .A3(_03417_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08087_ (.A1(_01123_),
    .A2(\register_file[30][27] ),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08088_ (.I(_01096_),
    .Z(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08089_ (.A1(_03420_),
    .A2(\register_file[31][27] ),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08090_ (.A1(_03419_),
    .A2(_01141_),
    .A3(_03421_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08091_ (.A1(_03418_),
    .A2(_03422_),
    .A3(_03340_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08092_ (.A1(_03415_),
    .A2(_03423_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08093_ (.A1(_03406_),
    .A2(_03424_),
    .A3(_03179_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08094_ (.A1(_03181_),
    .A2(\register_file[8][27] ),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08095_ (.A1(_03345_),
    .A2(\register_file[9][27] ),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08096_ (.A1(_03426_),
    .A2(_03427_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08097_ (.A1(_03428_),
    .A2(_03102_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08098_ (.A1(_03429_),
    .A2(_03104_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08099_ (.A1(_03350_),
    .A2(\register_file[11][27] ),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(_03352_),
    .A2(\register_file[10][27] ),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08101_ (.A1(_03431_),
    .A2(_03432_),
    .B(_03108_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08102_ (.A1(_03430_),
    .A2(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(_03356_),
    .A2(\register_file[12][27] ),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08104_ (.I(_01774_),
    .Z(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08105_ (.A1(_01048_),
    .A2(\register_file[13][27] ),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08106_ (.A1(_03435_),
    .A2(_03436_),
    .A3(_03437_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08107_ (.A1(_03274_),
    .A2(\register_file[14][27] ),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08108_ (.A1(_03276_),
    .A2(\register_file[15][27] ),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08109_ (.A1(_03439_),
    .A2(_03361_),
    .A3(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08110_ (.A1(_03438_),
    .A2(_03441_),
    .A3(_03279_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08111_ (.A1(_03434_),
    .A2(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08112_ (.A1(_03282_),
    .A2(\register_file[6][27] ),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08113_ (.I(\register_file[7][27] ),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08114_ (.A1(_03445_),
    .A2(_01167_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08115_ (.A1(_03444_),
    .A2(_03446_),
    .A3(_03369_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08116_ (.I(\register_file[4][27] ),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08117_ (.A1(_03203_),
    .A2(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08118_ (.I(\register_file[5][27] ),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08119_ (.A1(_03450_),
    .A2(_03374_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08120_ (.A1(_03449_),
    .A2(_03451_),
    .A3(_03376_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08121_ (.A1(_03447_),
    .A2(_03452_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08122_ (.A1(_03453_),
    .A2(_03210_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08123_ (.A1(_03380_),
    .A2(\register_file[2][27] ),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08124_ (.I(\register_file[3][27] ),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08125_ (.A1(_03456_),
    .A2(_03132_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08126_ (.A1(_03294_),
    .A2(_03455_),
    .A3(_03457_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08127_ (.I(_01005_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08128_ (.A1(_03459_),
    .A2(\register_file[1][27] ),
    .B(_01198_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08129_ (.A1(_03458_),
    .A2(_03460_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08130_ (.I(_03461_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08131_ (.A1(_03454_),
    .A2(_03462_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08132_ (.A1(_03443_),
    .A2(_03463_),
    .A3(_03303_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08133_ (.A1(_03425_),
    .A2(_03464_),
    .B(_03305_),
    .ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08134_ (.A1(_03306_),
    .A2(\register_file[24][28] ),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08135_ (.A1(_03222_),
    .A2(\register_file[25][28] ),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08136_ (.A1(_03465_),
    .A2(_03466_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08137_ (.A1(_03467_),
    .A2(_03225_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08138_ (.A1(_03468_),
    .A2(_01066_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08139_ (.A1(_01069_),
    .A2(\register_file[27][28] ),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08140_ (.A1(_03229_),
    .A2(\register_file[26][28] ),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08141_ (.A1(_03470_),
    .A2(_03471_),
    .B(_03231_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08142_ (.A1(_03469_),
    .A2(_03472_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08143_ (.A1(_01081_),
    .A2(\register_file[28][28] ),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08144_ (.A1(_03235_),
    .A2(\register_file[29][28] ),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08145_ (.A1(_03474_),
    .A2(_03150_),
    .A3(_03475_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08146_ (.A1(_03153_),
    .A2(\register_file[30][28] ),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08147_ (.A1(_03320_),
    .A2(\register_file[31][28] ),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08148_ (.A1(_03477_),
    .A2(_03155_),
    .A3(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08149_ (.A1(_03476_),
    .A2(_03479_),
    .A3(_01101_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08150_ (.A1(_03473_),
    .A2(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08151_ (.A1(_03243_),
    .A2(\register_file[16][28] ),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08152_ (.A1(_01111_),
    .A2(\register_file[17][28] ),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08153_ (.A1(_03482_),
    .A2(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08154_ (.A1(_03484_),
    .A2(_03163_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08155_ (.A1(_03485_),
    .A2(_01010_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08156_ (.A1(_01120_),
    .A2(\register_file[19][28] ),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08157_ (.A1(_01090_),
    .A2(\register_file[18][28] ),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08158_ (.A1(_03487_),
    .A2(_03488_),
    .B(_03168_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08159_ (.A1(_03486_),
    .A2(_03489_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08160_ (.A1(_01130_),
    .A2(\register_file[20][28] ),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08161_ (.A1(_01135_),
    .A2(\register_file[21][28] ),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08162_ (.A1(_03491_),
    .A2(_01133_),
    .A3(_03492_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08163_ (.A1(_01123_),
    .A2(\register_file[22][28] ),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08164_ (.A1(_03420_),
    .A2(\register_file[23][28] ),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08165_ (.A1(_03494_),
    .A2(_01141_),
    .A3(_03495_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08166_ (.A1(_03493_),
    .A2(_03496_),
    .A3(_03340_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08167_ (.A1(_03490_),
    .A2(_03497_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08168_ (.A1(_03481_),
    .A2(_03498_),
    .A3(_03179_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08169_ (.A1(_03181_),
    .A2(\register_file[8][28] ),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08170_ (.A1(_03345_),
    .A2(\register_file[9][28] ),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08171_ (.A1(_03500_),
    .A2(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08172_ (.A1(_03502_),
    .A2(_01186_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08173_ (.A1(_03503_),
    .A2(_01188_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08174_ (.A1(_03350_),
    .A2(\register_file[11][28] ),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08175_ (.A1(_03352_),
    .A2(\register_file[10][28] ),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08176_ (.A1(_03505_),
    .A2(_03506_),
    .B(_01025_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08177_ (.A1(_03504_),
    .A2(_03507_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08178_ (.A1(_03356_),
    .A2(\register_file[12][28] ),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08179_ (.A1(_01048_),
    .A2(\register_file[13][28] ),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08180_ (.A1(_03509_),
    .A2(_03436_),
    .A3(_03510_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08181_ (.A1(_03274_),
    .A2(\register_file[14][28] ),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08182_ (.A1(_03276_),
    .A2(\register_file[15][28] ),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08183_ (.A1(_03512_),
    .A2(_03361_),
    .A3(_03513_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08184_ (.A1(_03511_),
    .A2(_03514_),
    .A3(_03279_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08185_ (.A1(_03508_),
    .A2(_03515_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08186_ (.A1(_03282_),
    .A2(\register_file[6][28] ),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08187_ (.I(\register_file[7][28] ),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08188_ (.A1(_03518_),
    .A2(_01167_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08189_ (.A1(_03517_),
    .A2(_03519_),
    .A3(_03369_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08190_ (.I(\register_file[4][28] ),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08191_ (.A1(_03203_),
    .A2(_03521_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08192_ (.I(\register_file[5][28] ),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08193_ (.A1(_03523_),
    .A2(_03374_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08194_ (.A1(_03522_),
    .A2(_03524_),
    .A3(_03376_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08195_ (.A1(_03520_),
    .A2(_03525_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08196_ (.A1(_03526_),
    .A2(_03210_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08197_ (.A1(_03380_),
    .A2(\register_file[2][28] ),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08198_ (.I(\register_file[3][28] ),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08199_ (.A1(_03529_),
    .A2(_01156_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08200_ (.A1(_03294_),
    .A2(_03528_),
    .A3(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08201_ (.A1(_03459_),
    .A2(\register_file[1][28] ),
    .B(_01198_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08202_ (.A1(_03531_),
    .A2(_03532_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08203_ (.I(_03533_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08204_ (.A1(_03527_),
    .A2(_03534_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08205_ (.A1(_03516_),
    .A2(_03535_),
    .A3(_03303_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08206_ (.A1(_03499_),
    .A2(_03536_),
    .B(_03305_),
    .ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08207_ (.A1(_03306_),
    .A2(\register_file[16][29] ),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08208_ (.A1(_03222_),
    .A2(\register_file[17][29] ),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08209_ (.A1(_03537_),
    .A2(_03538_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08210_ (.A1(_03539_),
    .A2(_03225_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08211_ (.A1(_03540_),
    .A2(_02978_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08212_ (.A1(_01069_),
    .A2(\register_file[19][29] ),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08213_ (.A1(_03229_),
    .A2(\register_file[18][29] ),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08214_ (.A1(_03542_),
    .A2(_03543_),
    .B(_03231_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08215_ (.A1(_03541_),
    .A2(_03544_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08216_ (.A1(_01081_),
    .A2(\register_file[20][29] ),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08217_ (.A1(_03235_),
    .A2(\register_file[21][29] ),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08218_ (.A1(_03546_),
    .A2(_01084_),
    .A3(_03547_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08219_ (.A1(_01072_),
    .A2(\register_file[22][29] ),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08220_ (.A1(_03320_),
    .A2(\register_file[23][29] ),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08221_ (.A1(_03549_),
    .A2(_01094_),
    .A3(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08222_ (.A1(_03548_),
    .A2(_03551_),
    .A3(_01101_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08223_ (.A1(_03545_),
    .A2(_03552_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08224_ (.A1(_03243_),
    .A2(\register_file[24][29] ),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08225_ (.A1(_01111_),
    .A2(\register_file[25][29] ),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08226_ (.A1(_03554_),
    .A2(_03555_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08227_ (.A1(_03556_),
    .A2(_01115_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08228_ (.A1(_03557_),
    .A2(_01117_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08229_ (.A1(_01120_),
    .A2(\register_file[27][29] ),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08230_ (.A1(_01090_),
    .A2(\register_file[26][29] ),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08231_ (.A1(_03559_),
    .A2(_03560_),
    .B(_01126_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08232_ (.A1(_03558_),
    .A2(_03561_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08233_ (.A1(_01130_),
    .A2(\register_file[28][29] ),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08234_ (.A1(_01135_),
    .A2(\register_file[29][29] ),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08235_ (.A1(_03563_),
    .A2(_01133_),
    .A3(_03564_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08236_ (.A1(_01123_),
    .A2(\register_file[30][29] ),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08237_ (.A1(_03420_),
    .A2(\register_file[31][29] ),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08238_ (.A1(_03566_),
    .A2(_01141_),
    .A3(_03567_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08239_ (.A1(_03565_),
    .A2(_03568_),
    .A3(_03340_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08240_ (.A1(_03562_),
    .A2(_03569_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08241_ (.A1(_03553_),
    .A2(_03570_),
    .A3(_01505_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08242_ (.A1(_01030_),
    .A2(\register_file[8][29] ),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08243_ (.A1(_03345_),
    .A2(\register_file[9][29] ),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08244_ (.A1(_03572_),
    .A2(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08245_ (.A1(_03574_),
    .A2(_01186_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08246_ (.A1(_03575_),
    .A2(_01188_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08247_ (.A1(_03350_),
    .A2(\register_file[11][29] ),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08248_ (.A1(_03352_),
    .A2(\register_file[10][29] ),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08249_ (.A1(_03577_),
    .A2(_03578_),
    .B(_01025_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08250_ (.A1(_03576_),
    .A2(_03579_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08251_ (.A1(_03356_),
    .A2(\register_file[12][29] ),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08252_ (.A1(_01048_),
    .A2(\register_file[13][29] ),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08253_ (.A1(_03581_),
    .A2(_03436_),
    .A3(_03582_),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08254_ (.A1(_03274_),
    .A2(\register_file[14][29] ),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08255_ (.A1(_03276_),
    .A2(\register_file[15][29] ),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08256_ (.A1(_03584_),
    .A2(_03361_),
    .A3(_03585_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08257_ (.A1(_03583_),
    .A2(_03586_),
    .A3(_03279_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08258_ (.A1(_03580_),
    .A2(_03587_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08259_ (.A1(_03282_),
    .A2(\register_file[6][29] ),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08260_ (.I(\register_file[7][29] ),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08261_ (.A1(_03590_),
    .A2(_01167_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08262_ (.A1(_03589_),
    .A2(_03591_),
    .A3(_03369_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08263_ (.I(\register_file[4][29] ),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08264_ (.A1(_00995_),
    .A2(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08265_ (.I(\register_file[5][29] ),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08266_ (.A1(_03595_),
    .A2(_03374_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08267_ (.A1(_03594_),
    .A2(_03596_),
    .A3(_03376_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08268_ (.A1(_03592_),
    .A2(_03597_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08269_ (.A1(_03598_),
    .A2(_01052_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08270_ (.A1(_03380_),
    .A2(\register_file[2][29] ),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08271_ (.I(\register_file[3][29] ),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08272_ (.A1(_03601_),
    .A2(_01156_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08273_ (.A1(_03294_),
    .A2(_03600_),
    .A3(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08274_ (.A1(_03459_),
    .A2(\register_file[1][29] ),
    .B(_01198_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08275_ (.A1(_03603_),
    .A2(_03604_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08276_ (.I(_03605_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08277_ (.A1(_03599_),
    .A2(_03606_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08278_ (.A1(_03588_),
    .A2(_03607_),
    .A3(_03303_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08279_ (.A1(_03571_),
    .A2(_03608_),
    .B(_03305_),
    .ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08280_ (.A1(_03306_),
    .A2(\register_file[16][30] ),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08281_ (.A1(_01059_),
    .A2(\register_file[17][30] ),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08282_ (.A1(_03609_),
    .A2(_03610_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08283_ (.A1(_03611_),
    .A2(_01063_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08284_ (.A1(_03612_),
    .A2(_01490_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08285_ (.A1(_01069_),
    .A2(\register_file[19][30] ),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08286_ (.A1(_01043_),
    .A2(\register_file[18][30] ),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08287_ (.A1(_03614_),
    .A2(_03615_),
    .B(_01076_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08288_ (.A1(_03613_),
    .A2(_03616_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08289_ (.A1(_01081_),
    .A2(\register_file[20][30] ),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08290_ (.A1(_01086_),
    .A2(\register_file[21][30] ),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08291_ (.A1(_03618_),
    .A2(_01084_),
    .A3(_03619_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08292_ (.A1(_01072_),
    .A2(\register_file[22][30] ),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08293_ (.A1(_03320_),
    .A2(\register_file[23][30] ),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08294_ (.A1(_03621_),
    .A2(_01094_),
    .A3(_03622_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08295_ (.A1(_03620_),
    .A2(_03623_),
    .A3(_01101_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08296_ (.A1(_03617_),
    .A2(_03624_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08297_ (.A1(_01108_),
    .A2(\register_file[24][30] ),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08298_ (.A1(_01111_),
    .A2(\register_file[25][30] ),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08299_ (.A1(_03626_),
    .A2(_03627_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08300_ (.A1(_03628_),
    .A2(_01115_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08301_ (.A1(_03629_),
    .A2(_01117_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08302_ (.A1(_01120_),
    .A2(\register_file[27][30] ),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08303_ (.A1(_01090_),
    .A2(\register_file[26][30] ),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08304_ (.A1(_03631_),
    .A2(_03632_),
    .B(_01126_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08305_ (.A1(_03630_),
    .A2(_03633_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08306_ (.A1(_01130_),
    .A2(\register_file[28][30] ),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08307_ (.A1(_01135_),
    .A2(\register_file[29][30] ),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08308_ (.A1(_03635_),
    .A2(_01133_),
    .A3(_03636_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08309_ (.A1(_01123_),
    .A2(\register_file[30][30] ),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08310_ (.A1(_03420_),
    .A2(\register_file[31][30] ),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08311_ (.A1(_03638_),
    .A2(_01141_),
    .A3(_03639_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08312_ (.A1(_03637_),
    .A2(_03640_),
    .A3(_03340_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08313_ (.A1(_03634_),
    .A2(_03641_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08314_ (.A1(_03625_),
    .A2(_03642_),
    .A3(_01505_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08315_ (.A1(_01030_),
    .A2(\register_file[8][30] ),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08316_ (.A1(_03345_),
    .A2(\register_file[9][30] ),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08317_ (.A1(_03644_),
    .A2(_03645_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08318_ (.A1(_03646_),
    .A2(_01186_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08319_ (.A1(_03647_),
    .A2(_01188_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08320_ (.A1(_03350_),
    .A2(\register_file[11][30] ),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08321_ (.A1(_03352_),
    .A2(\register_file[10][30] ),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08322_ (.A1(_03649_),
    .A2(_03650_),
    .B(_01025_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08323_ (.A1(_03648_),
    .A2(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08324_ (.A1(_03356_),
    .A2(\register_file[12][30] ),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08325_ (.A1(_01048_),
    .A2(\register_file[13][30] ),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08326_ (.A1(_03653_),
    .A2(_03436_),
    .A3(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08327_ (.A1(_01162_),
    .A2(\register_file[14][30] ),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08328_ (.I(_01455_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08329_ (.A1(_03657_),
    .A2(\register_file[15][30] ),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08330_ (.A1(_03656_),
    .A2(_03361_),
    .A3(_03658_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08331_ (.A1(_03655_),
    .A2(_03659_),
    .A3(_01394_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08332_ (.A1(_03652_),
    .A2(_03660_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08333_ (.A1(_01179_),
    .A2(\register_file[6][30] ),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08334_ (.I(\register_file[7][30] ),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08335_ (.A1(_03663_),
    .A2(_01167_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08336_ (.A1(_03662_),
    .A2(_03664_),
    .A3(_03369_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08337_ (.I(\register_file[4][30] ),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08338_ (.A1(_00995_),
    .A2(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08339_ (.I(\register_file[5][30] ),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08340_ (.A1(_03668_),
    .A2(_03374_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08341_ (.A1(_03667_),
    .A2(_03669_),
    .A3(_03376_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08342_ (.A1(_03665_),
    .A2(_03670_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08343_ (.A1(_03671_),
    .A2(_01052_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08344_ (.A1(_03380_),
    .A2(\register_file[2][30] ),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08345_ (.I(\register_file[3][30] ),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08346_ (.A1(_03674_),
    .A2(_01156_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08347_ (.A1(_01176_),
    .A2(_03673_),
    .A3(_03675_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08348_ (.A1(_03459_),
    .A2(\register_file[1][30] ),
    .B(_01198_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08349_ (.A1(_03676_),
    .A2(_03677_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08350_ (.I(_03678_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08351_ (.A1(_03672_),
    .A2(_03679_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08352_ (.A1(_03661_),
    .A2(_03680_),
    .A3(_01194_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08353_ (.A1(_03643_),
    .A2(_03681_),
    .B(_01200_),
    .ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08354_ (.A1(_01179_),
    .A2(\register_file[6][31] ),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08355_ (.I(\register_file[7][31] ),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08356_ (.A1(_03683_),
    .A2(_01059_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08357_ (.A1(_03682_),
    .A2(_03684_),
    .A3(_01045_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08358_ (.I(\register_file[4][31] ),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08359_ (.A1(_00995_),
    .A2(_03686_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08360_ (.I(\register_file[5][31] ),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08361_ (.A1(_03688_),
    .A2(_01059_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08362_ (.A1(_03687_),
    .A2(_03689_),
    .A3(_01035_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08363_ (.A1(_03685_),
    .A2(_03690_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08364_ (.A1(_03691_),
    .A2(_01394_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08365_ (.A1(_00995_),
    .A2(\register_file[3][31] ),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08366_ (.A1(_03693_),
    .A2(_01025_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08367_ (.A1(_01182_),
    .A2(\register_file[2][31] ),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08368_ (.A1(_03459_),
    .A2(\register_file[1][31] ),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08369_ (.A1(_03694_),
    .A2(_03695_),
    .B(_03696_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08370_ (.A1(_03692_),
    .A2(_03697_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08371_ (.A1(_03698_),
    .A2(_01197_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08372_ (.A1(_03699_),
    .A2(_01011_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08373_ (.I(_01179_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08374_ (.A1(_03701_),
    .A2(\register_file[8][31] ),
    .Z(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08375_ (.I(\register_file[9][31] ),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08376_ (.A1(_03703_),
    .A2(_03420_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08377_ (.A1(_03702_),
    .A2(_03704_),
    .A3(_01170_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08378_ (.I(_01277_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08379_ (.A1(_03706_),
    .A2(\register_file[10][31] ),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08380_ (.I(\register_file[11][31] ),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08381_ (.A1(_03708_),
    .A2(_03657_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08382_ (.A1(_03707_),
    .A2(_03709_),
    .A3(_01159_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08383_ (.A1(_03705_),
    .A2(_03710_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08384_ (.A1(_03711_),
    .A2(_01022_),
    .B(_01011_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08385_ (.A1(_01031_),
    .A2(\register_file[12][31] ),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08386_ (.A1(_01015_),
    .A2(\register_file[13][31] ),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08387_ (.A1(_03713_),
    .A2(_01036_),
    .A3(_03714_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08388_ (.A1(_01031_),
    .A2(\register_file[14][31] ),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08389_ (.A1(_01015_),
    .A2(\register_file[15][31] ),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08390_ (.A1(_03716_),
    .A2(_01046_),
    .A3(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08391_ (.A1(_03715_),
    .A2(_03718_),
    .A3(_01173_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08392_ (.A1(_03712_),
    .A2(_03719_),
    .B(_01505_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08393_ (.A1(_03700_),
    .A2(_03720_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08394_ (.A1(_03701_),
    .A2(\register_file[30][31] ),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08395_ (.I(\register_file[31][31] ),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08396_ (.A1(_03723_),
    .A2(_01086_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08397_ (.A1(_03722_),
    .A2(_03724_),
    .A3(_01094_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08398_ (.A1(_03701_),
    .A2(\register_file[28][31] ),
    .Z(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08399_ (.I(\register_file[29][31] ),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08400_ (.A1(_03727_),
    .A2(_01097_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08401_ (.A1(_03726_),
    .A2(_03728_),
    .A3(_01170_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08402_ (.A1(_03725_),
    .A2(_03729_),
    .A3(_01101_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08403_ (.A1(_03701_),
    .A2(\register_file[24][31] ),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08404_ (.I(\register_file[25][31] ),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08405_ (.A1(_03732_),
    .A2(_01097_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08406_ (.A1(_03731_),
    .A2(_03733_),
    .A3(_01170_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08407_ (.A1(_03706_),
    .A2(\register_file[26][31] ),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08408_ (.I(\register_file[27][31] ),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08409_ (.A1(_03736_),
    .A2(_03657_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08410_ (.A1(_03735_),
    .A2(_03737_),
    .A3(_01159_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08411_ (.A1(_03734_),
    .A2(_03738_),
    .A3(_01022_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08412_ (.A1(_03730_),
    .A2(_03739_),
    .A3(_01468_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08413_ (.A1(_03701_),
    .A2(\register_file[16][31] ),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08414_ (.I(\register_file[17][31] ),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08415_ (.A1(_03742_),
    .A2(_01097_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08416_ (.A1(_03741_),
    .A2(_03743_),
    .A3(_03436_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08417_ (.A1(_03706_),
    .A2(\register_file[18][31] ),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08418_ (.I(\register_file[19][31] ),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08419_ (.A1(_03746_),
    .A2(_03657_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08420_ (.A1(_03745_),
    .A2(_03747_),
    .A3(_01159_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08421_ (.A1(_03744_),
    .A2(_03748_),
    .A3(_01022_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08422_ (.A1(_03706_),
    .A2(\register_file[22][31] ),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08423_ (.I(\register_file[23][31] ),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08424_ (.A1(_03751_),
    .A2(_03657_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08425_ (.A1(_03750_),
    .A2(_03752_),
    .A3(_01159_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08426_ (.A1(_03706_),
    .A2(\register_file[20][31] ),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08427_ (.I(\register_file[21][31] ),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08428_ (.A1(_03755_),
    .A2(_01182_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08429_ (.A1(_03754_),
    .A2(_03756_),
    .A3(_01170_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08430_ (.A1(_03753_),
    .A2(_03757_),
    .A3(_01394_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08431_ (.A1(_03749_),
    .A2(_03758_),
    .A3(_01011_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08432_ (.A1(_03740_),
    .A2(_03759_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08433_ (.A1(_03760_),
    .A2(_01105_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08434_ (.A1(_03721_),
    .A2(_03761_),
    .ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08435_ (.I(net2),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08436_ (.A1(_03762_),
    .A2(net1),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08437_ (.I(_03763_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08438_ (.I(_03764_),
    .Z(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08439_ (.I(_03765_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08440_ (.I(_03766_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08441_ (.A1(_03767_),
    .A2(\register_file[25][0] ),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08442_ (.A1(net1),
    .A2(net2),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08443_ (.I(_03769_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08444_ (.I(_03770_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08445_ (.I(_03771_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08446_ (.I(_03772_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08447_ (.A1(_03773_),
    .A2(\register_file[24][0] ),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08448_ (.A1(_03768_),
    .A2(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08449_ (.I(_03762_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08450_ (.A1(_03776_),
    .A2(net1),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08451_ (.I(_03777_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08452_ (.I(_03778_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08453_ (.I(_03779_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08454_ (.A1(_03780_),
    .A2(\register_file[26][0] ),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08455_ (.A1(net1),
    .A2(net2),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08456_ (.I(_03782_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08457_ (.I(_03783_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08458_ (.I(_03784_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08459_ (.I(_03785_),
    .Z(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08460_ (.A1(_03786_),
    .A2(\register_file[27][0] ),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08461_ (.A1(_03781_),
    .A2(_03787_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08462_ (.I(net5),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08463_ (.I(_03789_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08464_ (.I(net4),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08465_ (.I(_03791_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08466_ (.I(net3),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08467_ (.A1(_03790_),
    .A2(_03792_),
    .A3(_03793_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08468_ (.I(_03794_),
    .Z(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08469_ (.I(_03795_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08470_ (.A1(_03775_),
    .A2(_03788_),
    .B(_03796_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08471_ (.I(_03764_),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08472_ (.I(_03798_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08473_ (.I(_03799_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08474_ (.A1(_03800_),
    .A2(\register_file[29][0] ),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08475_ (.I(_03771_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08476_ (.I(_03802_),
    .Z(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08477_ (.A1(_03803_),
    .A2(\register_file[28][0] ),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08478_ (.A1(_03801_),
    .A2(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08479_ (.I(_03777_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08480_ (.I(_03806_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08481_ (.I(_03807_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08482_ (.A1(_03808_),
    .A2(\register_file[30][0] ),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08483_ (.I(_03784_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08484_ (.I(_03810_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08485_ (.A1(_03811_),
    .A2(\register_file[31][0] ),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08486_ (.A1(_03809_),
    .A2(_03812_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08487_ (.I(net3),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08488_ (.A1(_03790_),
    .A2(_03814_),
    .A3(_03792_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08489_ (.I(_03815_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08490_ (.I(_03816_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08491_ (.A1(_03805_),
    .A2(_03813_),
    .B(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08492_ (.A1(_03797_),
    .A2(_03818_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08493_ (.I(_03798_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08494_ (.I(_03820_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08495_ (.A1(_03821_),
    .A2(\register_file[21][0] ),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08496_ (.I(_03771_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08497_ (.I(_03823_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08498_ (.A1(_03824_),
    .A2(\register_file[20][0] ),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08499_ (.A1(_03822_),
    .A2(_03825_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08500_ (.I(_03778_),
    .Z(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08501_ (.I(_03827_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08502_ (.A1(_03828_),
    .A2(\register_file[22][0] ),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08503_ (.I(_03783_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08504_ (.I(_03830_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08505_ (.I(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08506_ (.A1(_03832_),
    .A2(\register_file[23][0] ),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08507_ (.A1(_03829_),
    .A2(_03833_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08508_ (.A1(_03792_),
    .A2(net5),
    .A3(_03793_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08509_ (.I(_03835_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08510_ (.I(_03836_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08511_ (.I(_03837_),
    .Z(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08512_ (.A1(_03826_),
    .A2(_03834_),
    .B(_03838_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08513_ (.I(_03798_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08514_ (.I(_03840_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08515_ (.A1(_03841_),
    .A2(\register_file[17][0] ),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08516_ (.I(_03770_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08517_ (.I(_03843_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08518_ (.A1(_03844_),
    .A2(\register_file[16][0] ),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08519_ (.A1(_03842_),
    .A2(_03845_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08520_ (.I(_03806_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08521_ (.I(_03847_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08522_ (.A1(_03848_),
    .A2(\register_file[18][0] ),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08523_ (.I(_03784_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08524_ (.I(_03850_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08525_ (.A1(_03851_),
    .A2(\register_file[19][0] ),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08526_ (.A1(_03849_),
    .A2(_03852_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08527_ (.A1(_03790_),
    .A2(_03793_),
    .A3(net4),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08528_ (.I(_03854_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08529_ (.I(_03855_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08530_ (.A1(_03846_),
    .A2(_03853_),
    .B(_03856_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08531_ (.A1(_03839_),
    .A2(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08532_ (.A1(_03819_),
    .A2(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08533_ (.I(_03798_),
    .Z(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08534_ (.I(_03860_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08535_ (.A1(_03861_),
    .A2(\register_file[13][0] ),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08536_ (.I(_03771_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08537_ (.I(_03863_),
    .Z(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08538_ (.A1(_03864_),
    .A2(\register_file[12][0] ),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08539_ (.A1(_03862_),
    .A2(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08540_ (.I(_03806_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08541_ (.I(_03867_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08542_ (.A1(_03868_),
    .A2(\register_file[14][0] ),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08543_ (.I(_03784_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08544_ (.I(_03870_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08545_ (.A1(_03871_),
    .A2(\register_file[15][0] ),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08546_ (.A1(_03869_),
    .A2(_03872_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08547_ (.A1(_03790_),
    .A2(_03793_),
    .A3(net4),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08548_ (.I(_03874_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08549_ (.I(_03875_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08550_ (.I(_03876_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08551_ (.A1(_03866_),
    .A2(_03873_),
    .B(_03877_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08552_ (.I(_03764_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08553_ (.I(_03879_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08554_ (.A1(_03880_),
    .A2(\register_file[9][0] ),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08555_ (.I(_03770_),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08556_ (.I(_03882_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08557_ (.A1(_03883_),
    .A2(\register_file[8][0] ),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08558_ (.A1(_03881_),
    .A2(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08559_ (.I(_03777_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08560_ (.I(_03886_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08561_ (.A1(_03887_),
    .A2(\register_file[10][0] ),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08562_ (.I(_03783_),
    .Z(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08563_ (.I(_03889_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08564_ (.A1(_03890_),
    .A2(\register_file[11][0] ),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08565_ (.A1(_03888_),
    .A2(_03891_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08566_ (.A1(_03792_),
    .A2(net5),
    .A3(_03793_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08567_ (.I(_03893_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08568_ (.A1(_03885_),
    .A2(_03892_),
    .B(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08569_ (.A1(_03878_),
    .A2(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08570_ (.I(_03764_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08571_ (.I(_03897_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08572_ (.A1(_03898_),
    .A2(\register_file[5][0] ),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08573_ (.I(_03770_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08574_ (.I(_03900_),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08575_ (.A1(_03901_),
    .A2(\register_file[4][0] ),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08576_ (.A1(_03899_),
    .A2(_03902_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08577_ (.I(_03806_),
    .Z(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08578_ (.I(_03904_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08579_ (.A1(_03905_),
    .A2(\register_file[6][0] ),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08580_ (.I(_03784_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08581_ (.I(_03907_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08582_ (.A1(_03908_),
    .A2(\register_file[7][0] ),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08583_ (.A1(_03906_),
    .A2(_03909_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08584_ (.A1(_03789_),
    .A2(_03791_),
    .A3(net3),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08585_ (.I(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08586_ (.I(_03912_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08587_ (.I(_03913_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08588_ (.A1(_03903_),
    .A2(_03910_),
    .B(_03914_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08589_ (.I(_03806_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08590_ (.I(_03916_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08591_ (.A1(_03917_),
    .A2(\register_file[2][0] ),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08592_ (.I(_03830_),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08593_ (.I(_03919_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08594_ (.A1(_03920_),
    .A2(\register_file[3][0] ),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08595_ (.I(_03776_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08596_ (.I(_03922_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08597_ (.A1(_03923_),
    .A2(\register_file[1][0] ),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08598_ (.A1(_03918_),
    .A2(_03921_),
    .A3(_03924_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08599_ (.A1(_03790_),
    .A2(_03814_),
    .A3(_03792_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08600_ (.I(_03926_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08601_ (.I(_03927_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08602_ (.I(_03928_),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08603_ (.A1(_03925_),
    .A2(_03929_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08604_ (.A1(_03915_),
    .A2(_03930_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08605_ (.A1(_03896_),
    .A2(_03931_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08606_ (.I(_03772_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08607_ (.A1(_03928_),
    .A2(_03933_),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08608_ (.I(_03934_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08609_ (.I(_03935_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08610_ (.A1(_03859_),
    .A2(_03932_),
    .B(_03936_),
    .ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08611_ (.A1(_03767_),
    .A2(\register_file[29][1] ),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08612_ (.A1(_03773_),
    .A2(\register_file[28][1] ),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08613_ (.A1(_03937_),
    .A2(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08614_ (.A1(_03780_),
    .A2(\register_file[30][1] ),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08615_ (.A1(_03786_),
    .A2(\register_file[31][1] ),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08616_ (.A1(_03940_),
    .A2(_03941_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08617_ (.I(_03816_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08618_ (.A1(_03939_),
    .A2(_03942_),
    .B(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08619_ (.A1(_03800_),
    .A2(\register_file[25][1] ),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08620_ (.A1(_03803_),
    .A2(\register_file[24][1] ),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08621_ (.A1(_03945_),
    .A2(_03946_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08622_ (.A1(_03808_),
    .A2(\register_file[26][1] ),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08623_ (.A1(_03811_),
    .A2(\register_file[27][1] ),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08624_ (.A1(_03948_),
    .A2(_03949_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08625_ (.A1(_03947_),
    .A2(_03950_),
    .B(_03796_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08626_ (.A1(_03944_),
    .A2(_03951_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08627_ (.A1(_03821_),
    .A2(\register_file[5][1] ),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08628_ (.A1(_03824_),
    .A2(\register_file[4][1] ),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08629_ (.A1(_03953_),
    .A2(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08630_ (.I(_03827_),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08631_ (.A1(_03956_),
    .A2(\register_file[6][1] ),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08632_ (.I(_03831_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08633_ (.A1(_03958_),
    .A2(\register_file[7][1] ),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08634_ (.A1(_03957_),
    .A2(_03959_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08635_ (.I(_03912_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08636_ (.I(_03961_),
    .Z(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08637_ (.A1(_03955_),
    .A2(_03960_),
    .B(_03962_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08638_ (.I(_03798_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08639_ (.I(_03964_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08640_ (.A1(_03965_),
    .A2(\register_file[17][1] ),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08641_ (.I(_03843_),
    .Z(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08642_ (.A1(_03967_),
    .A2(\register_file[16][1] ),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08643_ (.A1(_03966_),
    .A2(_03968_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08644_ (.A1(_03848_),
    .A2(\register_file[18][1] ),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08645_ (.A1(_03851_),
    .A2(\register_file[19][1] ),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08646_ (.A1(_03970_),
    .A2(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08647_ (.A1(_03969_),
    .A2(_03972_),
    .B(_03856_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08648_ (.A1(_03963_),
    .A2(_03973_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08649_ (.A1(_03952_),
    .A2(_03974_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08650_ (.A1(_03861_),
    .A2(\register_file[13][1] ),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08651_ (.A1(_03864_),
    .A2(\register_file[12][1] ),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08652_ (.A1(_03976_),
    .A2(_03977_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08653_ (.A1(_03868_),
    .A2(\register_file[14][1] ),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08654_ (.A1(_03871_),
    .A2(\register_file[15][1] ),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08655_ (.A1(_03979_),
    .A2(_03980_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08656_ (.A1(_03978_),
    .A2(_03981_),
    .B(_03877_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08657_ (.A1(_03880_),
    .A2(\register_file[21][1] ),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08658_ (.A1(_03883_),
    .A2(\register_file[20][1] ),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08659_ (.A1(_03983_),
    .A2(_03984_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08660_ (.I(_03886_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08661_ (.A1(_03986_),
    .A2(\register_file[22][1] ),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08662_ (.I(_03889_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08663_ (.A1(_03988_),
    .A2(\register_file[23][1] ),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08664_ (.A1(_03987_),
    .A2(_03989_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08665_ (.I(_03836_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08666_ (.I(_03991_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08667_ (.A1(_03985_),
    .A2(_03990_),
    .B(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08668_ (.A1(_03982_),
    .A2(_03993_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08669_ (.A1(_03898_),
    .A2(\register_file[9][1] ),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08670_ (.A1(_03901_),
    .A2(\register_file[8][1] ),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08671_ (.A1(_03995_),
    .A2(_03996_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08672_ (.A1(_03905_),
    .A2(\register_file[10][1] ),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08673_ (.A1(_03908_),
    .A2(\register_file[11][1] ),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08674_ (.A1(_03998_),
    .A2(_03999_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08675_ (.I(_03893_),
    .Z(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08676_ (.I(_04001_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08677_ (.A1(_03997_),
    .A2(_04000_),
    .B(_04002_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08678_ (.A1(_03917_),
    .A2(\register_file[2][1] ),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08679_ (.A1(_03920_),
    .A2(\register_file[3][1] ),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08680_ (.A1(_03923_),
    .A2(\register_file[1][1] ),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08681_ (.A1(_04004_),
    .A2(_04005_),
    .A3(_04006_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08682_ (.A1(_04007_),
    .A2(_03929_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08683_ (.A1(_04003_),
    .A2(_04008_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08684_ (.A1(_03994_),
    .A2(_04009_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08685_ (.A1(_03975_),
    .A2(_04010_),
    .B(_03936_),
    .ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08686_ (.A1(_03767_),
    .A2(\register_file[17][2] ),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08687_ (.A1(_03773_),
    .A2(\register_file[16][2] ),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08688_ (.A1(_04011_),
    .A2(_04012_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08689_ (.A1(_03780_),
    .A2(\register_file[18][2] ),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08690_ (.A1(_03786_),
    .A2(\register_file[19][2] ),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08691_ (.A1(_04014_),
    .A2(_04015_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08692_ (.I(_03854_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08693_ (.I(_04017_),
    .Z(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08694_ (.A1(_04013_),
    .A2(_04016_),
    .B(_04018_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08695_ (.A1(_03800_),
    .A2(\register_file[21][2] ),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08696_ (.A1(_03803_),
    .A2(\register_file[20][2] ),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08697_ (.A1(_04020_),
    .A2(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08698_ (.A1(_03808_),
    .A2(\register_file[22][2] ),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08699_ (.A1(_03811_),
    .A2(\register_file[23][2] ),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08700_ (.A1(_04023_),
    .A2(_04024_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08701_ (.I(_03837_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08702_ (.A1(_04022_),
    .A2(_04025_),
    .B(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08703_ (.A1(_04019_),
    .A2(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08704_ (.I(_03820_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08705_ (.A1(_04029_),
    .A2(\register_file[9][2] ),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08706_ (.I(_03823_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08707_ (.A1(_04031_),
    .A2(\register_file[8][2] ),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08708_ (.A1(_04030_),
    .A2(_04032_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08709_ (.A1(_03956_),
    .A2(\register_file[10][2] ),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08710_ (.A1(_03958_),
    .A2(\register_file[11][2] ),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08711_ (.A1(_04034_),
    .A2(_04035_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08712_ (.I(_03894_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08713_ (.A1(_04033_),
    .A2(_04036_),
    .B(_04037_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08714_ (.A1(_03965_),
    .A2(\register_file[13][2] ),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08715_ (.A1(_03967_),
    .A2(\register_file[12][2] ),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08716_ (.A1(_04039_),
    .A2(_04040_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08717_ (.A1(_03848_),
    .A2(\register_file[14][2] ),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08718_ (.A1(_03851_),
    .A2(\register_file[15][2] ),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08719_ (.A1(_04042_),
    .A2(_04043_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08720_ (.I(_03876_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08721_ (.A1(_04041_),
    .A2(_04044_),
    .B(_04045_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08722_ (.A1(_04038_),
    .A2(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08723_ (.A1(_04028_),
    .A2(_04047_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08724_ (.A1(_03861_),
    .A2(\register_file[5][2] ),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08725_ (.A1(_03864_),
    .A2(\register_file[4][2] ),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08726_ (.A1(_04049_),
    .A2(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08727_ (.I(_03867_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08728_ (.A1(_04052_),
    .A2(\register_file[6][2] ),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08729_ (.I(_03870_),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08730_ (.A1(_04054_),
    .A2(\register_file[7][2] ),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08731_ (.A1(_04053_),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08732_ (.I(_03913_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08733_ (.A1(_04051_),
    .A2(_04056_),
    .B(_04057_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08734_ (.I(_03879_),
    .Z(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08735_ (.A1(_04059_),
    .A2(\register_file[25][2] ),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08736_ (.I(_03882_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08737_ (.A1(_04061_),
    .A2(\register_file[24][2] ),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08738_ (.A1(_04060_),
    .A2(_04062_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08739_ (.A1(_03986_),
    .A2(\register_file[26][2] ),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08740_ (.A1(_03988_),
    .A2(\register_file[27][2] ),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08741_ (.A1(_04064_),
    .A2(_04065_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08742_ (.I(_03794_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08743_ (.I(_04067_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08744_ (.A1(_04063_),
    .A2(_04066_),
    .B(_04068_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08745_ (.A1(_04058_),
    .A2(_04069_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08746_ (.A1(_03898_),
    .A2(\register_file[29][2] ),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08747_ (.A1(_03901_),
    .A2(\register_file[28][2] ),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08748_ (.A1(_04071_),
    .A2(_04072_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08749_ (.A1(_03905_),
    .A2(\register_file[30][2] ),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08750_ (.A1(_03908_),
    .A2(\register_file[31][2] ),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08751_ (.A1(_04074_),
    .A2(_04075_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08752_ (.I(_03815_),
    .Z(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08753_ (.I(_04077_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08754_ (.A1(_04073_),
    .A2(_04076_),
    .B(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08755_ (.A1(_03917_),
    .A2(\register_file[2][2] ),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08756_ (.A1(_03920_),
    .A2(\register_file[3][2] ),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08757_ (.A1(_03923_),
    .A2(\register_file[1][2] ),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08758_ (.A1(_04080_),
    .A2(_04081_),
    .A3(_04082_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08759_ (.A1(_04083_),
    .A2(_03929_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08760_ (.A1(_04079_),
    .A2(_04084_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08761_ (.A1(_04070_),
    .A2(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08762_ (.A1(_04048_),
    .A2(_04086_),
    .B(_03936_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08763_ (.A1(_03767_),
    .A2(\register_file[13][3] ),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08764_ (.A1(_03773_),
    .A2(\register_file[12][3] ),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08765_ (.A1(_04087_),
    .A2(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08766_ (.I(_03779_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08767_ (.A1(_04090_),
    .A2(\register_file[14][3] ),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08768_ (.A1(_03786_),
    .A2(\register_file[15][3] ),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08769_ (.A1(_04091_),
    .A2(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08770_ (.I(_03876_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08771_ (.A1(_04089_),
    .A2(_04093_),
    .B(_04094_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08772_ (.A1(_03800_),
    .A2(\register_file[17][3] ),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08773_ (.A1(_03803_),
    .A2(\register_file[16][3] ),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08774_ (.A1(_04096_),
    .A2(_04097_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08775_ (.A1(_03808_),
    .A2(\register_file[18][3] ),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08776_ (.A1(_03811_),
    .A2(\register_file[19][3] ),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08777_ (.A1(_04099_),
    .A2(_04100_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08778_ (.I(_04017_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08779_ (.A1(_04098_),
    .A2(_04101_),
    .B(_04102_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08780_ (.A1(_04095_),
    .A2(_04103_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08781_ (.A1(_04029_),
    .A2(\register_file[21][3] ),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08782_ (.A1(_04031_),
    .A2(\register_file[20][3] ),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08783_ (.A1(_04105_),
    .A2(_04106_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08784_ (.A1(_03956_),
    .A2(\register_file[22][3] ),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08785_ (.A1(_03958_),
    .A2(\register_file[23][3] ),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08786_ (.A1(_04108_),
    .A2(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08787_ (.A1(_04107_),
    .A2(_04110_),
    .B(_03838_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08788_ (.A1(_03965_),
    .A2(\register_file[9][3] ),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08789_ (.A1(_03967_),
    .A2(\register_file[8][3] ),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08790_ (.A1(_04112_),
    .A2(_04113_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08791_ (.A1(_03848_),
    .A2(\register_file[10][3] ),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08792_ (.A1(_03851_),
    .A2(\register_file[11][3] ),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08793_ (.A1(_04115_),
    .A2(_04116_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08794_ (.I(_04001_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08795_ (.A1(_04114_),
    .A2(_04117_),
    .B(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08796_ (.A1(_04111_),
    .A2(_04119_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08797_ (.A1(_04104_),
    .A2(_04120_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08798_ (.I(_03860_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08799_ (.A1(_04122_),
    .A2(\register_file[25][3] ),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08800_ (.I(_03771_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08801_ (.I(_04124_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08802_ (.A1(_04125_),
    .A2(\register_file[24][3] ),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08803_ (.A1(_04123_),
    .A2(_04126_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08804_ (.A1(_04052_),
    .A2(\register_file[26][3] ),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08805_ (.A1(_04054_),
    .A2(\register_file[27][3] ),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08806_ (.A1(_04128_),
    .A2(_04129_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08807_ (.I(_03795_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08808_ (.A1(_04127_),
    .A2(_04130_),
    .B(_04131_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08809_ (.A1(_04059_),
    .A2(\register_file[29][3] ),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08810_ (.A1(_04061_),
    .A2(\register_file[28][3] ),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08811_ (.A1(_04133_),
    .A2(_04134_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08812_ (.A1(_03986_),
    .A2(\register_file[30][3] ),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08813_ (.A1(_03988_),
    .A2(\register_file[31][3] ),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08814_ (.A1(_04136_),
    .A2(_04137_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08815_ (.I(_04077_),
    .Z(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08816_ (.A1(_04135_),
    .A2(_04138_),
    .B(_04139_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08817_ (.A1(_04132_),
    .A2(_04140_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08818_ (.A1(_03898_),
    .A2(\register_file[5][3] ),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08819_ (.A1(_03901_),
    .A2(\register_file[4][3] ),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08820_ (.A1(_04142_),
    .A2(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08821_ (.I(_03777_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08822_ (.I(_04145_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08823_ (.A1(_04146_),
    .A2(\register_file[6][3] ),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08824_ (.I(_03783_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08825_ (.I(_04148_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08826_ (.A1(_04149_),
    .A2(\register_file[7][3] ),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08827_ (.A1(_04147_),
    .A2(_04150_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08828_ (.A1(_04144_),
    .A2(_04151_),
    .B(_03914_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08829_ (.A1(_03917_),
    .A2(\register_file[2][3] ),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08830_ (.I(_03919_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08831_ (.A1(_04154_),
    .A2(\register_file[3][3] ),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08832_ (.A1(_03923_),
    .A2(\register_file[1][3] ),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08833_ (.A1(_04153_),
    .A2(_04155_),
    .A3(_04156_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08834_ (.A1(_04157_),
    .A2(_03929_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08835_ (.A1(_04152_),
    .A2(_04158_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08836_ (.A1(_04141_),
    .A2(_04159_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08837_ (.A1(_04121_),
    .A2(_04160_),
    .B(_03936_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08838_ (.A1(_03933_),
    .A2(\register_file[4][4] ),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08839_ (.A1(_01534_),
    .A2(_03763_),
    .B(_04161_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08840_ (.A1(_04090_),
    .A2(\register_file[6][4] ),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08841_ (.A1(_03786_),
    .A2(\register_file[7][4] ),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08842_ (.A1(_04163_),
    .A2(_04164_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08843_ (.A1(_04162_),
    .A2(_04165_),
    .B(_03962_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08844_ (.A1(_03800_),
    .A2(\register_file[17][4] ),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08845_ (.A1(_03803_),
    .A2(\register_file[16][4] ),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08846_ (.A1(_04167_),
    .A2(_04168_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08847_ (.I(_03807_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08848_ (.A1(_04170_),
    .A2(\register_file[18][4] ),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08849_ (.I(_03810_),
    .Z(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08850_ (.A1(_04172_),
    .A2(\register_file[19][4] ),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08851_ (.A1(_04171_),
    .A2(_04173_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08852_ (.A1(_04169_),
    .A2(_04174_),
    .B(_04102_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08853_ (.A1(_04166_),
    .A2(_04175_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08854_ (.A1(_04029_),
    .A2(\register_file[29][4] ),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08855_ (.A1(_04031_),
    .A2(\register_file[28][4] ),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08856_ (.A1(_04177_),
    .A2(_04178_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08857_ (.A1(_03956_),
    .A2(\register_file[30][4] ),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08858_ (.A1(_03958_),
    .A2(\register_file[31][4] ),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08859_ (.A1(_04180_),
    .A2(_04181_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08860_ (.I(_03816_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08861_ (.A1(_04179_),
    .A2(_04182_),
    .B(_04183_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08862_ (.A1(_03965_),
    .A2(\register_file[25][4] ),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08863_ (.A1(_03967_),
    .A2(\register_file[24][4] ),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08864_ (.A1(_04185_),
    .A2(_04186_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08865_ (.A1(_03848_),
    .A2(\register_file[26][4] ),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08866_ (.A1(_03851_),
    .A2(\register_file[27][4] ),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08867_ (.A1(_04188_),
    .A2(_04189_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08868_ (.I(_04067_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08869_ (.A1(_04187_),
    .A2(_04190_),
    .B(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08870_ (.A1(_04184_),
    .A2(_04192_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08871_ (.A1(_04176_),
    .A2(_04193_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08872_ (.A1(_04122_),
    .A2(\register_file[9][4] ),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08873_ (.A1(_04125_),
    .A2(\register_file[8][4] ),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08874_ (.A1(_04195_),
    .A2(_04196_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08875_ (.A1(_04052_),
    .A2(\register_file[10][4] ),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08876_ (.A1(_04054_),
    .A2(\register_file[11][4] ),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08877_ (.A1(_04198_),
    .A2(_04199_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08878_ (.I(_03894_),
    .Z(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08879_ (.A1(_04197_),
    .A2(_04200_),
    .B(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08880_ (.A1(_04059_),
    .A2(\register_file[21][4] ),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08881_ (.A1(_04061_),
    .A2(\register_file[20][4] ),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08882_ (.A1(_04203_),
    .A2(_04204_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08883_ (.A1(_03986_),
    .A2(\register_file[22][4] ),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08884_ (.A1(_03988_),
    .A2(\register_file[23][4] ),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08885_ (.A1(_04206_),
    .A2(_04207_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08886_ (.A1(_04205_),
    .A2(_04208_),
    .B(_03992_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08887_ (.A1(_04202_),
    .A2(_04209_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08888_ (.I(_03897_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08889_ (.A1(_04211_),
    .A2(\register_file[13][4] ),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08890_ (.I(_03900_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08891_ (.A1(_04213_),
    .A2(\register_file[12][4] ),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08892_ (.A1(_04212_),
    .A2(_04214_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08893_ (.A1(_04146_),
    .A2(\register_file[14][4] ),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08894_ (.A1(_04149_),
    .A2(\register_file[15][4] ),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08895_ (.A1(_04216_),
    .A2(_04217_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08896_ (.I(_03875_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08897_ (.I(_04219_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08898_ (.A1(_04215_),
    .A2(_04218_),
    .B(_04220_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08899_ (.A1(_03917_),
    .A2(\register_file[2][4] ),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08900_ (.A1(_04154_),
    .A2(\register_file[3][4] ),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08901_ (.A1(_03923_),
    .A2(\register_file[1][4] ),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08902_ (.A1(_04222_),
    .A2(_04223_),
    .A3(_04224_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08903_ (.A1(_04225_),
    .A2(_03929_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08904_ (.A1(_04221_),
    .A2(_04226_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08905_ (.A1(_04210_),
    .A2(_04227_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08906_ (.A1(_04194_),
    .A2(_04228_),
    .B(_03936_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08907_ (.A1(_03767_),
    .A2(\register_file[9][5] ),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08908_ (.A1(_03773_),
    .A2(\register_file[8][5] ),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08909_ (.A1(_04229_),
    .A2(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08910_ (.A1(_04090_),
    .A2(\register_file[10][5] ),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08911_ (.I(_03785_),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(_04233_),
    .A2(\register_file[11][5] ),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08913_ (.A1(_04232_),
    .A2(_04234_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08914_ (.A1(_04231_),
    .A2(_04235_),
    .B(_04037_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08915_ (.I(_03799_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08916_ (.A1(_04237_),
    .A2(\register_file[17][5] ),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08917_ (.I(_03802_),
    .Z(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(_04239_),
    .A2(\register_file[16][5] ),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08919_ (.A1(_04238_),
    .A2(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08920_ (.A1(_04170_),
    .A2(\register_file[18][5] ),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08921_ (.A1(_04172_),
    .A2(\register_file[19][5] ),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08922_ (.A1(_04242_),
    .A2(_04243_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08923_ (.A1(_04241_),
    .A2(_04244_),
    .B(_04102_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08924_ (.A1(_04236_),
    .A2(_04245_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08925_ (.A1(_04029_),
    .A2(\register_file[13][5] ),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08926_ (.A1(_04031_),
    .A2(\register_file[12][5] ),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08927_ (.A1(_04247_),
    .A2(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08928_ (.A1(_03956_),
    .A2(\register_file[14][5] ),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08929_ (.A1(_03958_),
    .A2(\register_file[15][5] ),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08930_ (.A1(_04250_),
    .A2(_04251_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08931_ (.A1(_04249_),
    .A2(_04252_),
    .B(_03877_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08932_ (.A1(_03965_),
    .A2(\register_file[21][5] ),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08933_ (.A1(_03967_),
    .A2(\register_file[20][5] ),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08934_ (.A1(_04254_),
    .A2(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08935_ (.I(_03847_),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08936_ (.A1(_04257_),
    .A2(\register_file[22][5] ),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08937_ (.I(_03850_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08938_ (.A1(_04259_),
    .A2(\register_file[23][5] ),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08939_ (.A1(_04258_),
    .A2(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08940_ (.I(_03837_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08941_ (.A1(_04256_),
    .A2(_04261_),
    .B(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08942_ (.A1(_04253_),
    .A2(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08943_ (.A1(_04246_),
    .A2(_04264_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08944_ (.A1(_04122_),
    .A2(\register_file[29][5] ),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08945_ (.A1(_04125_),
    .A2(\register_file[28][5] ),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08946_ (.A1(_04266_),
    .A2(_04267_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08947_ (.A1(_04052_),
    .A2(\register_file[30][5] ),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08948_ (.A1(_04054_),
    .A2(\register_file[31][5] ),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08949_ (.A1(_04269_),
    .A2(_04270_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08950_ (.A1(_04268_),
    .A2(_04271_),
    .B(_03817_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08951_ (.A1(_04059_),
    .A2(\register_file[25][5] ),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08952_ (.A1(_04061_),
    .A2(\register_file[24][5] ),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08953_ (.A1(_04273_),
    .A2(_04274_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08954_ (.A1(_03986_),
    .A2(\register_file[26][5] ),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08955_ (.A1(_03988_),
    .A2(\register_file[27][5] ),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08956_ (.A1(_04276_),
    .A2(_04277_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08957_ (.A1(_04275_),
    .A2(_04278_),
    .B(_04068_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08958_ (.A1(_04272_),
    .A2(_04279_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08959_ (.A1(_04211_),
    .A2(\register_file[5][5] ),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08960_ (.A1(_04213_),
    .A2(\register_file[4][5] ),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08961_ (.A1(_04281_),
    .A2(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08962_ (.A1(_04146_),
    .A2(\register_file[6][5] ),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08963_ (.A1(_04149_),
    .A2(\register_file[7][5] ),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08964_ (.A1(_04284_),
    .A2(_04285_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08965_ (.A1(_04283_),
    .A2(_04286_),
    .B(_03914_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08966_ (.I(_03916_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08967_ (.A1(_04288_),
    .A2(\register_file[2][5] ),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08968_ (.A1(_04154_),
    .A2(\register_file[3][5] ),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08969_ (.I(_03922_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08970_ (.A1(_04291_),
    .A2(\register_file[1][5] ),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08971_ (.A1(_04289_),
    .A2(_04290_),
    .A3(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08972_ (.I(_03928_),
    .Z(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08973_ (.A1(_04293_),
    .A2(_04294_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08974_ (.A1(_04287_),
    .A2(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08975_ (.A1(_04280_),
    .A2(_04296_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08976_ (.I(_03935_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08977_ (.A1(_04265_),
    .A2(_04297_),
    .B(_04298_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08978_ (.A1(_03933_),
    .A2(\register_file[4][6] ),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08979_ (.A1(_01706_),
    .A2(_03763_),
    .B(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08980_ (.A1(_04090_),
    .A2(\register_file[6][6] ),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08981_ (.A1(_04233_),
    .A2(\register_file[7][6] ),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08982_ (.A1(_04301_),
    .A2(_04302_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08983_ (.A1(_04300_),
    .A2(_04303_),
    .B(_03962_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08984_ (.A1(_04237_),
    .A2(\register_file[29][6] ),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08985_ (.A1(_04239_),
    .A2(\register_file[28][6] ),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08986_ (.A1(_04305_),
    .A2(_04306_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08987_ (.A1(_04170_),
    .A2(\register_file[30][6] ),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08988_ (.A1(_04172_),
    .A2(\register_file[31][6] ),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08989_ (.A1(_04308_),
    .A2(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08990_ (.A1(_04307_),
    .A2(_04310_),
    .B(_03817_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08991_ (.A1(_04304_),
    .A2(_04311_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08992_ (.A1(_04029_),
    .A2(\register_file[17][6] ),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08993_ (.A1(_04031_),
    .A2(\register_file[16][6] ),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08994_ (.A1(_04313_),
    .A2(_04314_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08995_ (.I(_03778_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08996_ (.I(_04316_),
    .Z(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08997_ (.A1(_04317_),
    .A2(\register_file[18][6] ),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08998_ (.I(_03830_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08999_ (.I(_04319_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09000_ (.A1(_04320_),
    .A2(\register_file[19][6] ),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09001_ (.A1(_04318_),
    .A2(_04321_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09002_ (.I(_04017_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09003_ (.A1(_04315_),
    .A2(_04322_),
    .B(_04323_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09004_ (.I(_03964_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09005_ (.A1(_04325_),
    .A2(\register_file[21][6] ),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09006_ (.I(_03843_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09007_ (.A1(_04327_),
    .A2(\register_file[20][6] ),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09008_ (.A1(_04326_),
    .A2(_04328_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09009_ (.A1(_04257_),
    .A2(\register_file[22][6] ),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09010_ (.A1(_04259_),
    .A2(\register_file[23][6] ),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09011_ (.A1(_04330_),
    .A2(_04331_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09012_ (.A1(_04329_),
    .A2(_04332_),
    .B(_04262_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09013_ (.A1(_04324_),
    .A2(_04333_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09014_ (.A1(_04312_),
    .A2(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09015_ (.A1(_04122_),
    .A2(\register_file[9][6] ),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09016_ (.A1(_04125_),
    .A2(\register_file[8][6] ),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09017_ (.A1(_04336_),
    .A2(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09018_ (.A1(_04052_),
    .A2(\register_file[10][6] ),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09019_ (.A1(_04054_),
    .A2(\register_file[11][6] ),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09020_ (.A1(_04339_),
    .A2(_04340_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09021_ (.A1(_04338_),
    .A2(_04341_),
    .B(_04201_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09022_ (.A1(_04059_),
    .A2(\register_file[25][6] ),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09023_ (.A1(_04061_),
    .A2(\register_file[24][6] ),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09024_ (.A1(_04343_),
    .A2(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09025_ (.I(_03886_),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09026_ (.A1(_04346_),
    .A2(\register_file[26][6] ),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09027_ (.I(_03889_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09028_ (.A1(_04348_),
    .A2(\register_file[27][6] ),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09029_ (.A1(_04347_),
    .A2(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09030_ (.A1(_04345_),
    .A2(_04350_),
    .B(_04068_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09031_ (.A1(_04342_),
    .A2(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09032_ (.A1(_04211_),
    .A2(\register_file[13][6] ),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(_04213_),
    .A2(\register_file[12][6] ),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09034_ (.A1(_04353_),
    .A2(_04354_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09035_ (.A1(_04146_),
    .A2(\register_file[14][6] ),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09036_ (.A1(_04149_),
    .A2(\register_file[15][6] ),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09037_ (.A1(_04356_),
    .A2(_04357_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09038_ (.A1(_04355_),
    .A2(_04358_),
    .B(_04220_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09039_ (.A1(_04288_),
    .A2(\register_file[2][6] ),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09040_ (.A1(_04154_),
    .A2(\register_file[3][6] ),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09041_ (.A1(_04291_),
    .A2(\register_file[1][6] ),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09042_ (.A1(_04360_),
    .A2(_04361_),
    .A3(_04362_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09043_ (.A1(_04363_),
    .A2(_04294_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09044_ (.A1(_04359_),
    .A2(_04364_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09045_ (.A1(_04352_),
    .A2(_04365_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09046_ (.A1(_04335_),
    .A2(_04366_),
    .B(_04298_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09047_ (.I(_03766_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09048_ (.A1(_04367_),
    .A2(\register_file[13][7] ),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09049_ (.I(_03772_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09050_ (.A1(_04369_),
    .A2(\register_file[12][7] ),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09051_ (.A1(_04368_),
    .A2(_04370_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09052_ (.A1(_04090_),
    .A2(\register_file[14][7] ),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09053_ (.A1(_04233_),
    .A2(\register_file[15][7] ),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09054_ (.A1(_04372_),
    .A2(_04373_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09055_ (.A1(_04371_),
    .A2(_04374_),
    .B(_04094_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09056_ (.A1(_04237_),
    .A2(\register_file[25][7] ),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09057_ (.A1(_04239_),
    .A2(\register_file[24][7] ),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09058_ (.A1(_04376_),
    .A2(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09059_ (.A1(_04170_),
    .A2(\register_file[26][7] ),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09060_ (.A1(_04172_),
    .A2(\register_file[27][7] ),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09061_ (.A1(_04379_),
    .A2(_04380_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09062_ (.I(_03795_),
    .Z(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09063_ (.A1(_04378_),
    .A2(_04381_),
    .B(_04382_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09064_ (.A1(_04375_),
    .A2(_04383_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09065_ (.I(_03820_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09066_ (.A1(_04385_),
    .A2(\register_file[17][7] ),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09067_ (.I(_03823_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09068_ (.A1(_04387_),
    .A2(\register_file[16][7] ),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09069_ (.A1(_04386_),
    .A2(_04388_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09070_ (.A1(_04317_),
    .A2(\register_file[18][7] ),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09071_ (.A1(_04320_),
    .A2(\register_file[19][7] ),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09072_ (.A1(_04390_),
    .A2(_04391_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09073_ (.A1(_04389_),
    .A2(_04392_),
    .B(_04323_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09074_ (.A1(_04325_),
    .A2(\register_file[21][7] ),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09075_ (.A1(_04327_),
    .A2(\register_file[20][7] ),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09076_ (.A1(_04394_),
    .A2(_04395_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09077_ (.A1(_04257_),
    .A2(\register_file[22][7] ),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09078_ (.A1(_04259_),
    .A2(\register_file[23][7] ),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09079_ (.A1(_04397_),
    .A2(_04398_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09080_ (.I(_03991_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09081_ (.A1(_04396_),
    .A2(_04399_),
    .B(_04400_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09082_ (.A1(_04393_),
    .A2(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09083_ (.A1(_04384_),
    .A2(_04402_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09084_ (.A1(_04122_),
    .A2(\register_file[9][7] ),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09085_ (.A1(_04125_),
    .A2(\register_file[8][7] ),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09086_ (.A1(_04404_),
    .A2(_04405_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09087_ (.I(_03867_),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09088_ (.A1(_04407_),
    .A2(\register_file[10][7] ),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09089_ (.I(_03870_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09090_ (.A1(_04409_),
    .A2(\register_file[11][7] ),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09091_ (.A1(_04408_),
    .A2(_04410_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09092_ (.A1(_04406_),
    .A2(_04411_),
    .B(_04201_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09093_ (.I(_03879_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09094_ (.A1(_04413_),
    .A2(\register_file[5][7] ),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09095_ (.I(_03770_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09096_ (.I(_04415_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09097_ (.A1(_04416_),
    .A2(\register_file[4][7] ),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09098_ (.A1(_04414_),
    .A2(_04417_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09099_ (.A1(_04346_),
    .A2(\register_file[6][7] ),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09100_ (.A1(_04348_),
    .A2(\register_file[7][7] ),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09101_ (.A1(_04419_),
    .A2(_04420_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09102_ (.A1(_04418_),
    .A2(_04421_),
    .B(_03961_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09103_ (.A1(_04412_),
    .A2(_04422_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09104_ (.A1(_04211_),
    .A2(\register_file[29][7] ),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09105_ (.A1(_04213_),
    .A2(\register_file[28][7] ),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09106_ (.A1(_04424_),
    .A2(_04425_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09107_ (.A1(_04146_),
    .A2(\register_file[30][7] ),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09108_ (.A1(_04149_),
    .A2(\register_file[31][7] ),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09109_ (.A1(_04427_),
    .A2(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09110_ (.A1(_04426_),
    .A2(_04429_),
    .B(_04078_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09111_ (.A1(_04288_),
    .A2(\register_file[2][7] ),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09112_ (.A1(_04154_),
    .A2(\register_file[3][7] ),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09113_ (.A1(_04291_),
    .A2(\register_file[1][7] ),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09114_ (.A1(_04431_),
    .A2(_04432_),
    .A3(_04433_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09115_ (.A1(_04434_),
    .A2(_04294_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09116_ (.A1(_04430_),
    .A2(_04435_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09117_ (.A1(_04423_),
    .A2(_04436_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09118_ (.A1(_04403_),
    .A2(_04437_),
    .B(_04298_),
    .ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09119_ (.A1(_04367_),
    .A2(\register_file[29][8] ),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09120_ (.A1(_04369_),
    .A2(\register_file[28][8] ),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09121_ (.A1(_04438_),
    .A2(_04439_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09122_ (.I(_03779_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09123_ (.A1(_04441_),
    .A2(\register_file[30][8] ),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09124_ (.A1(_04233_),
    .A2(\register_file[31][8] ),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09125_ (.A1(_04442_),
    .A2(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09126_ (.A1(_04440_),
    .A2(_04444_),
    .B(_03943_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09127_ (.A1(_04237_),
    .A2(\register_file[17][8] ),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09128_ (.A1(_04239_),
    .A2(\register_file[16][8] ),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09129_ (.A1(_04446_),
    .A2(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09130_ (.A1(_04170_),
    .A2(\register_file[18][8] ),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09131_ (.A1(_04172_),
    .A2(\register_file[19][8] ),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09132_ (.A1(_04449_),
    .A2(_04450_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09133_ (.I(_03855_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09134_ (.A1(_04448_),
    .A2(_04451_),
    .B(_04452_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09135_ (.A1(_04445_),
    .A2(_04453_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09136_ (.A1(_04385_),
    .A2(\register_file[5][8] ),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09137_ (.A1(_04387_),
    .A2(\register_file[4][8] ),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09138_ (.A1(_04455_),
    .A2(_04456_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09139_ (.A1(_04317_),
    .A2(\register_file[6][8] ),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09140_ (.A1(_04320_),
    .A2(\register_file[7][8] ),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09141_ (.A1(_04458_),
    .A2(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09142_ (.A1(_04457_),
    .A2(_04460_),
    .B(_03962_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09143_ (.A1(_04325_),
    .A2(\register_file[21][8] ),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09144_ (.A1(_04327_),
    .A2(\register_file[20][8] ),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09145_ (.A1(_04462_),
    .A2(_04463_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09146_ (.A1(_04257_),
    .A2(\register_file[22][8] ),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09147_ (.A1(_04259_),
    .A2(\register_file[23][8] ),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09148_ (.A1(_04465_),
    .A2(_04466_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09149_ (.A1(_04464_),
    .A2(_04467_),
    .B(_04400_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09150_ (.A1(_04461_),
    .A2(_04468_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09151_ (.A1(_04454_),
    .A2(_04469_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09152_ (.I(_03840_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09153_ (.A1(_04471_),
    .A2(\register_file[9][8] ),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09154_ (.I(_04124_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09155_ (.A1(_04473_),
    .A2(\register_file[8][8] ),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09156_ (.A1(_04472_),
    .A2(_04474_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09157_ (.A1(_04407_),
    .A2(\register_file[10][8] ),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09158_ (.A1(_04409_),
    .A2(\register_file[11][8] ),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09159_ (.A1(_04476_),
    .A2(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09160_ (.A1(_04475_),
    .A2(_04478_),
    .B(_04201_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09161_ (.A1(_04413_),
    .A2(\register_file[25][8] ),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09162_ (.A1(_04416_),
    .A2(\register_file[24][8] ),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09163_ (.A1(_04480_),
    .A2(_04481_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09164_ (.A1(_04346_),
    .A2(\register_file[26][8] ),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09165_ (.A1(_04348_),
    .A2(\register_file[27][8] ),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09166_ (.A1(_04483_),
    .A2(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09167_ (.I(_04067_),
    .Z(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09168_ (.A1(_04482_),
    .A2(_04485_),
    .B(_04486_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09169_ (.A1(_04479_),
    .A2(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09170_ (.A1(_04211_),
    .A2(\register_file[13][8] ),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09171_ (.A1(_04213_),
    .A2(\register_file[12][8] ),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09172_ (.A1(_04489_),
    .A2(_04490_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09173_ (.I(_04145_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09174_ (.A1(_04492_),
    .A2(\register_file[14][8] ),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09175_ (.I(_04148_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09176_ (.A1(_04494_),
    .A2(\register_file[15][8] ),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09177_ (.A1(_04493_),
    .A2(_04495_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09178_ (.A1(_04491_),
    .A2(_04496_),
    .B(_04220_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09179_ (.A1(_04288_),
    .A2(\register_file[2][8] ),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09180_ (.I(_03919_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09181_ (.A1(_04499_),
    .A2(\register_file[3][8] ),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09182_ (.A1(_04291_),
    .A2(\register_file[1][8] ),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09183_ (.A1(_04498_),
    .A2(_04500_),
    .A3(_04501_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09184_ (.A1(_04502_),
    .A2(_04294_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09185_ (.A1(_04497_),
    .A2(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09186_ (.A1(_04488_),
    .A2(_04504_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09187_ (.A1(_04470_),
    .A2(_04505_),
    .B(_04298_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09188_ (.A1(_04367_),
    .A2(\register_file[13][9] ),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09189_ (.A1(_04369_),
    .A2(\register_file[12][9] ),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09190_ (.A1(_04506_),
    .A2(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09191_ (.A1(_04441_),
    .A2(\register_file[14][9] ),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09192_ (.A1(_04233_),
    .A2(\register_file[15][9] ),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(_04509_),
    .A2(_04510_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09194_ (.A1(_04508_),
    .A2(_04511_),
    .B(_04094_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(_04237_),
    .A2(\register_file[25][9] ),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09196_ (.A1(_04239_),
    .A2(\register_file[24][9] ),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09197_ (.A1(_04513_),
    .A2(_04514_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09198_ (.I(_03807_),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09199_ (.A1(_04516_),
    .A2(\register_file[26][9] ),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09200_ (.I(_03810_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09201_ (.A1(_04518_),
    .A2(\register_file[27][9] ),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09202_ (.A1(_04517_),
    .A2(_04519_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09203_ (.A1(_04515_),
    .A2(_04520_),
    .B(_04382_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09204_ (.A1(_04512_),
    .A2(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09205_ (.A1(_04385_),
    .A2(\register_file[5][9] ),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09206_ (.A1(_04387_),
    .A2(\register_file[4][9] ),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09207_ (.A1(_04523_),
    .A2(_04524_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09208_ (.A1(_04317_),
    .A2(\register_file[6][9] ),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09209_ (.A1(_04320_),
    .A2(\register_file[7][9] ),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09210_ (.A1(_04526_),
    .A2(_04527_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09211_ (.I(_03961_),
    .Z(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09212_ (.A1(_04525_),
    .A2(_04528_),
    .B(_04529_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09213_ (.A1(_04325_),
    .A2(\register_file[21][9] ),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09214_ (.A1(_04327_),
    .A2(\register_file[20][9] ),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(_04531_),
    .A2(_04532_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09216_ (.A1(_04257_),
    .A2(\register_file[22][9] ),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09217_ (.A1(_04259_),
    .A2(\register_file[23][9] ),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09218_ (.A1(_04534_),
    .A2(_04535_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09219_ (.A1(_04533_),
    .A2(_04536_),
    .B(_04400_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09220_ (.A1(_04530_),
    .A2(_04537_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09221_ (.A1(_04522_),
    .A2(_04538_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09222_ (.A1(_04471_),
    .A2(\register_file[9][9] ),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09223_ (.A1(_04473_),
    .A2(\register_file[8][9] ),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09224_ (.A1(_04540_),
    .A2(_04541_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09225_ (.A1(_04407_),
    .A2(\register_file[10][9] ),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09226_ (.A1(_04409_),
    .A2(\register_file[11][9] ),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09227_ (.A1(_04543_),
    .A2(_04544_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09228_ (.A1(_04542_),
    .A2(_04545_),
    .B(_04118_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09229_ (.A1(_04413_),
    .A2(\register_file[17][9] ),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09230_ (.A1(_04416_),
    .A2(\register_file[16][9] ),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09231_ (.A1(_04547_),
    .A2(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09232_ (.A1(_04346_),
    .A2(\register_file[18][9] ),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(_04348_),
    .A2(\register_file[19][9] ),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09234_ (.A1(_04550_),
    .A2(_04551_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09235_ (.I(_03855_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09236_ (.A1(_04549_),
    .A2(_04552_),
    .B(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09237_ (.A1(_04546_),
    .A2(_04554_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09238_ (.I(_03897_),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09239_ (.A1(_04556_),
    .A2(\register_file[29][9] ),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09240_ (.I(_03900_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09241_ (.A1(_04558_),
    .A2(\register_file[28][9] ),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09242_ (.A1(_04557_),
    .A2(_04559_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09243_ (.A1(_04492_),
    .A2(\register_file[30][9] ),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09244_ (.A1(_04494_),
    .A2(\register_file[31][9] ),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09245_ (.A1(_04561_),
    .A2(_04562_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09246_ (.A1(_04560_),
    .A2(_04563_),
    .B(_04078_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09247_ (.A1(_04288_),
    .A2(\register_file[2][9] ),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09248_ (.A1(_04499_),
    .A2(\register_file[3][9] ),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09249_ (.A1(_04291_),
    .A2(\register_file[1][9] ),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09250_ (.A1(_04565_),
    .A2(_04566_),
    .A3(_04567_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09251_ (.A1(_04568_),
    .A2(_04294_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09252_ (.A1(_04564_),
    .A2(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09253_ (.A1(_04555_),
    .A2(_04570_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09254_ (.A1(_04539_),
    .A2(_04571_),
    .B(_04298_),
    .ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09255_ (.A1(_04367_),
    .A2(\register_file[29][10] ),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09256_ (.A1(_04369_),
    .A2(\register_file[28][10] ),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09257_ (.A1(_04572_),
    .A2(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09258_ (.A1(_04441_),
    .A2(\register_file[30][10] ),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09259_ (.I(_03785_),
    .Z(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(_04576_),
    .A2(\register_file[31][10] ),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09261_ (.A1(_04575_),
    .A2(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09262_ (.A1(_04574_),
    .A2(_04578_),
    .B(_03943_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09263_ (.I(_03799_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09264_ (.A1(_04580_),
    .A2(\register_file[21][10] ),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09265_ (.I(_03863_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09266_ (.A1(_04582_),
    .A2(\register_file[20][10] ),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09267_ (.A1(_04581_),
    .A2(_04583_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09268_ (.A1(_04516_),
    .A2(\register_file[22][10] ),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09269_ (.A1(_04518_),
    .A2(\register_file[23][10] ),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09270_ (.A1(_04585_),
    .A2(_04586_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09271_ (.A1(_04584_),
    .A2(_04587_),
    .B(_04026_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09272_ (.A1(_04579_),
    .A2(_04588_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09273_ (.A1(_04385_),
    .A2(\register_file[5][10] ),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09274_ (.A1(_04387_),
    .A2(\register_file[4][10] ),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09275_ (.A1(_04590_),
    .A2(_04591_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09276_ (.A1(_04317_),
    .A2(\register_file[6][10] ),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09277_ (.A1(_04320_),
    .A2(\register_file[7][10] ),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(_04593_),
    .A2(_04594_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09279_ (.A1(_04592_),
    .A2(_04595_),
    .B(_04529_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09280_ (.A1(_04325_),
    .A2(\register_file[17][10] ),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09281_ (.A1(_04327_),
    .A2(\register_file[16][10] ),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09282_ (.A1(_04597_),
    .A2(_04598_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09283_ (.I(_03904_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09284_ (.A1(_04600_),
    .A2(\register_file[18][10] ),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09285_ (.I(_03907_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09286_ (.A1(_04602_),
    .A2(\register_file[19][10] ),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09287_ (.A1(_04601_),
    .A2(_04603_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09288_ (.A1(_04599_),
    .A2(_04604_),
    .B(_03856_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09289_ (.A1(_04596_),
    .A2(_04605_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09290_ (.A1(_04589_),
    .A2(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09291_ (.A1(_04471_),
    .A2(\register_file[13][10] ),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09292_ (.A1(_04473_),
    .A2(\register_file[12][10] ),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09293_ (.A1(_04608_),
    .A2(_04609_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09294_ (.A1(_04407_),
    .A2(\register_file[14][10] ),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09295_ (.A1(_04409_),
    .A2(\register_file[15][10] ),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(_04611_),
    .A2(_04612_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09297_ (.A1(_04610_),
    .A2(_04613_),
    .B(_04045_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09298_ (.A1(_04413_),
    .A2(\register_file[25][10] ),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09299_ (.A1(_04416_),
    .A2(\register_file[24][10] ),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09300_ (.A1(_04615_),
    .A2(_04616_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09301_ (.A1(_04346_),
    .A2(\register_file[26][10] ),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09302_ (.A1(_04348_),
    .A2(\register_file[27][10] ),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09303_ (.A1(_04618_),
    .A2(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09304_ (.A1(_04617_),
    .A2(_04620_),
    .B(_04486_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09305_ (.A1(_04614_),
    .A2(_04621_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09306_ (.A1(_04556_),
    .A2(\register_file[9][10] ),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09307_ (.A1(_04558_),
    .A2(\register_file[8][10] ),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09308_ (.A1(_04623_),
    .A2(_04624_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09309_ (.A1(_04492_),
    .A2(\register_file[10][10] ),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09310_ (.A1(_04494_),
    .A2(\register_file[11][10] ),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09311_ (.A1(_04626_),
    .A2(_04627_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09312_ (.A1(_04625_),
    .A2(_04628_),
    .B(_04002_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09313_ (.I(_03916_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09314_ (.A1(_04630_),
    .A2(\register_file[2][10] ),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(_04499_),
    .A2(\register_file[3][10] ),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09316_ (.I(_03922_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09317_ (.A1(_04633_),
    .A2(\register_file[1][10] ),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09318_ (.A1(_04631_),
    .A2(_04632_),
    .A3(_04634_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09319_ (.I(_03927_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09320_ (.I(_04636_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09321_ (.A1(_04635_),
    .A2(_04637_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09322_ (.A1(_04629_),
    .A2(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09323_ (.A1(_04622_),
    .A2(_04639_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09324_ (.I(_03935_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09325_ (.A1(_04607_),
    .A2(_04640_),
    .B(_04641_),
    .ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09326_ (.A1(_04367_),
    .A2(\register_file[25][11] ),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09327_ (.A1(_04369_),
    .A2(\register_file[24][11] ),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(_04642_),
    .A2(_04643_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09329_ (.A1(_04441_),
    .A2(\register_file[26][11] ),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09330_ (.A1(_04576_),
    .A2(\register_file[27][11] ),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09331_ (.A1(_04645_),
    .A2(_04646_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09332_ (.A1(_04644_),
    .A2(_04647_),
    .B(_03796_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09333_ (.A1(_04580_),
    .A2(\register_file[5][11] ),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09334_ (.A1(_04582_),
    .A2(\register_file[4][11] ),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09335_ (.A1(_04649_),
    .A2(_04650_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09336_ (.A1(_04516_),
    .A2(\register_file[6][11] ),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09337_ (.A1(_04518_),
    .A2(\register_file[7][11] ),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09338_ (.A1(_04652_),
    .A2(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09339_ (.I(_03961_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09340_ (.A1(_04651_),
    .A2(_04654_),
    .B(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09341_ (.A1(_04648_),
    .A2(_04656_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09342_ (.A1(_04385_),
    .A2(\register_file[21][11] ),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09343_ (.A1(_04387_),
    .A2(\register_file[20][11] ),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09344_ (.A1(_04658_),
    .A2(_04659_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09345_ (.I(_04316_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09346_ (.A1(_04661_),
    .A2(\register_file[22][11] ),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09347_ (.I(_04319_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09348_ (.A1(_04663_),
    .A2(\register_file[23][11] ),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09349_ (.A1(_04662_),
    .A2(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09350_ (.A1(_04660_),
    .A2(_04665_),
    .B(_03838_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09351_ (.I(_03964_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09352_ (.A1(_04667_),
    .A2(\register_file[29][11] ),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09353_ (.I(_03843_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09354_ (.A1(_04669_),
    .A2(\register_file[28][11] ),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09355_ (.A1(_04668_),
    .A2(_04670_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09356_ (.A1(_04600_),
    .A2(\register_file[30][11] ),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09357_ (.A1(_04602_),
    .A2(\register_file[31][11] ),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09358_ (.A1(_04672_),
    .A2(_04673_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09359_ (.I(_04077_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09360_ (.A1(_04671_),
    .A2(_04674_),
    .B(_04675_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09361_ (.A1(_04666_),
    .A2(_04676_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09362_ (.A1(_04657_),
    .A2(_04677_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09363_ (.A1(_04471_),
    .A2(\register_file[13][11] ),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09364_ (.A1(_04473_),
    .A2(\register_file[12][11] ),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09365_ (.A1(_04679_),
    .A2(_04680_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09366_ (.A1(_04407_),
    .A2(\register_file[14][11] ),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09367_ (.A1(_04409_),
    .A2(\register_file[15][11] ),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09368_ (.A1(_04682_),
    .A2(_04683_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09369_ (.A1(_04681_),
    .A2(_04684_),
    .B(_04045_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09370_ (.A1(_04413_),
    .A2(\register_file[9][11] ),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09371_ (.A1(_04416_),
    .A2(\register_file[8][11] ),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09372_ (.A1(_04686_),
    .A2(_04687_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09373_ (.I(_03886_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09374_ (.A1(_04689_),
    .A2(\register_file[10][11] ),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09375_ (.I(_03889_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09376_ (.A1(_04691_),
    .A2(\register_file[11][11] ),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09377_ (.A1(_04690_),
    .A2(_04692_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09378_ (.A1(_04688_),
    .A2(_04693_),
    .B(_03894_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09379_ (.A1(_04685_),
    .A2(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09380_ (.A1(_04556_),
    .A2(\register_file[17][11] ),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09381_ (.A1(_04558_),
    .A2(\register_file[16][11] ),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09382_ (.A1(_04696_),
    .A2(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09383_ (.A1(_04492_),
    .A2(\register_file[18][11] ),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09384_ (.A1(_04494_),
    .A2(\register_file[19][11] ),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09385_ (.A1(_04699_),
    .A2(_04700_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09386_ (.A1(_04698_),
    .A2(_04701_),
    .B(_04553_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09387_ (.A1(_04630_),
    .A2(\register_file[2][11] ),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09388_ (.A1(_04499_),
    .A2(\register_file[3][11] ),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09389_ (.A1(_04633_),
    .A2(\register_file[1][11] ),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09390_ (.A1(_04703_),
    .A2(_04704_),
    .A3(_04705_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09391_ (.A1(_04706_),
    .A2(_04637_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09392_ (.A1(_04702_),
    .A2(_04707_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09393_ (.A1(_04695_),
    .A2(_04708_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09394_ (.A1(_04678_),
    .A2(_04709_),
    .B(_04641_),
    .ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09395_ (.I(_03766_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09396_ (.A1(_04710_),
    .A2(\register_file[17][12] ),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09397_ (.I(_03772_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09398_ (.A1(_04712_),
    .A2(\register_file[16][12] ),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09399_ (.A1(_04711_),
    .A2(_04713_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09400_ (.A1(_04441_),
    .A2(\register_file[18][12] ),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09401_ (.A1(_04576_),
    .A2(\register_file[19][12] ),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09402_ (.A1(_04715_),
    .A2(_04716_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09403_ (.A1(_04714_),
    .A2(_04717_),
    .B(_04018_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09404_ (.A1(_04580_),
    .A2(\register_file[29][12] ),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09405_ (.A1(_04582_),
    .A2(\register_file[28][12] ),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09406_ (.A1(_04719_),
    .A2(_04720_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09407_ (.A1(_04516_),
    .A2(\register_file[30][12] ),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09408_ (.A1(_04518_),
    .A2(\register_file[31][12] ),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09409_ (.A1(_04722_),
    .A2(_04723_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09410_ (.A1(_04721_),
    .A2(_04724_),
    .B(_03817_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09411_ (.A1(_04718_),
    .A2(_04725_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09412_ (.I(_03820_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09413_ (.A1(_04727_),
    .A2(\register_file[5][12] ),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09414_ (.I(_03823_),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09415_ (.A1(_04729_),
    .A2(\register_file[4][12] ),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09416_ (.A1(_04728_),
    .A2(_04730_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09417_ (.A1(_04661_),
    .A2(\register_file[6][12] ),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09418_ (.A1(_04663_),
    .A2(\register_file[7][12] ),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09419_ (.A1(_04732_),
    .A2(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09420_ (.A1(_04731_),
    .A2(_04734_),
    .B(_04529_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09421_ (.A1(_04667_),
    .A2(\register_file[21][12] ),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09422_ (.A1(_04669_),
    .A2(\register_file[20][12] ),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09423_ (.A1(_04736_),
    .A2(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09424_ (.A1(_04600_),
    .A2(\register_file[22][12] ),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09425_ (.A1(_04602_),
    .A2(\register_file[23][12] ),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09426_ (.A1(_04739_),
    .A2(_04740_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09427_ (.A1(_04738_),
    .A2(_04741_),
    .B(_04400_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09428_ (.A1(_04735_),
    .A2(_04742_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09429_ (.A1(_04726_),
    .A2(_04743_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09430_ (.A1(_04471_),
    .A2(\register_file[9][12] ),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09431_ (.A1(_04473_),
    .A2(\register_file[8][12] ),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09432_ (.A1(_04745_),
    .A2(_04746_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09433_ (.I(_03867_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09434_ (.A1(_04748_),
    .A2(\register_file[10][12] ),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09435_ (.I(_03870_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09436_ (.A1(_04750_),
    .A2(\register_file[11][12] ),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09437_ (.A1(_04749_),
    .A2(_04751_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09438_ (.A1(_04747_),
    .A2(_04752_),
    .B(_04118_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09439_ (.I(_03765_),
    .Z(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09440_ (.A1(_04754_),
    .A2(\register_file[25][12] ),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09441_ (.I(_04415_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09442_ (.A1(_04756_),
    .A2(\register_file[24][12] ),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09443_ (.A1(_04755_),
    .A2(_04757_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09444_ (.A1(_04689_),
    .A2(\register_file[26][12] ),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09445_ (.A1(_04691_),
    .A2(\register_file[27][12] ),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09446_ (.A1(_04759_),
    .A2(_04760_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09447_ (.A1(_04758_),
    .A2(_04761_),
    .B(_04486_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09448_ (.A1(_04753_),
    .A2(_04762_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09449_ (.A1(_04556_),
    .A2(\register_file[13][12] ),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09450_ (.A1(_04558_),
    .A2(\register_file[12][12] ),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09451_ (.A1(_04764_),
    .A2(_04765_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09452_ (.A1(_04492_),
    .A2(\register_file[14][12] ),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09453_ (.A1(_04494_),
    .A2(\register_file[15][12] ),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09454_ (.A1(_04767_),
    .A2(_04768_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09455_ (.A1(_04766_),
    .A2(_04769_),
    .B(_04220_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09456_ (.A1(_04630_),
    .A2(\register_file[2][12] ),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09457_ (.A1(_04499_),
    .A2(\register_file[3][12] ),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09458_ (.A1(_04633_),
    .A2(\register_file[1][12] ),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09459_ (.A1(_04771_),
    .A2(_04772_),
    .A3(_04773_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(_04774_),
    .A2(_04637_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09461_ (.A1(_04770_),
    .A2(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09462_ (.A1(_04763_),
    .A2(_04776_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09463_ (.A1(_04744_),
    .A2(_04777_),
    .B(_04641_),
    .ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09464_ (.A1(_04710_),
    .A2(\register_file[13][13] ),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09465_ (.A1(_04712_),
    .A2(\register_file[12][13] ),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09466_ (.A1(_04778_),
    .A2(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09467_ (.I(_03827_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09468_ (.A1(_04781_),
    .A2(\register_file[14][13] ),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09469_ (.A1(_04576_),
    .A2(\register_file[15][13] ),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09470_ (.A1(_04782_),
    .A2(_04783_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09471_ (.A1(_04780_),
    .A2(_04784_),
    .B(_04094_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09472_ (.A1(_04580_),
    .A2(\register_file[25][13] ),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09473_ (.A1(_04582_),
    .A2(\register_file[24][13] ),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09474_ (.A1(_04786_),
    .A2(_04787_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09475_ (.A1(_04516_),
    .A2(\register_file[26][13] ),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09476_ (.A1(_04518_),
    .A2(\register_file[27][13] ),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09477_ (.A1(_04789_),
    .A2(_04790_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09478_ (.A1(_04788_),
    .A2(_04791_),
    .B(_04382_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09479_ (.A1(_04785_),
    .A2(_04792_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09480_ (.A1(_04727_),
    .A2(\register_file[17][13] ),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09481_ (.A1(_04729_),
    .A2(\register_file[16][13] ),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09482_ (.A1(_04794_),
    .A2(_04795_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09483_ (.A1(_04661_),
    .A2(\register_file[18][13] ),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(_04663_),
    .A2(\register_file[19][13] ),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09485_ (.A1(_04797_),
    .A2(_04798_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09486_ (.A1(_04796_),
    .A2(_04799_),
    .B(_04102_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09487_ (.A1(_04667_),
    .A2(\register_file[21][13] ),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09488_ (.A1(_04669_),
    .A2(\register_file[20][13] ),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09489_ (.A1(_04801_),
    .A2(_04802_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(_04600_),
    .A2(\register_file[22][13] ),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09491_ (.A1(_04602_),
    .A2(\register_file[23][13] ),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09492_ (.A1(_04804_),
    .A2(_04805_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09493_ (.A1(_04803_),
    .A2(_04806_),
    .B(_04400_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09494_ (.A1(_04800_),
    .A2(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09495_ (.A1(_04793_),
    .A2(_04808_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09496_ (.I(_03840_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09497_ (.A1(_04810_),
    .A2(\register_file[5][13] ),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09498_ (.I(_04124_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09499_ (.A1(_04812_),
    .A2(\register_file[4][13] ),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09500_ (.A1(_04811_),
    .A2(_04813_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09501_ (.A1(_04748_),
    .A2(\register_file[6][13] ),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09502_ (.A1(_04750_),
    .A2(\register_file[7][13] ),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09503_ (.A1(_04815_),
    .A2(_04816_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09504_ (.A1(_04814_),
    .A2(_04817_),
    .B(_04057_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09505_ (.A1(_04754_),
    .A2(\register_file[29][13] ),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09506_ (.A1(_04756_),
    .A2(\register_file[28][13] ),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09507_ (.A1(_04819_),
    .A2(_04820_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09508_ (.A1(_04689_),
    .A2(\register_file[30][13] ),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09509_ (.A1(_04691_),
    .A2(\register_file[31][13] ),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09510_ (.A1(_04822_),
    .A2(_04823_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09511_ (.A1(_04821_),
    .A2(_04824_),
    .B(_04139_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09512_ (.A1(_04818_),
    .A2(_04825_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09513_ (.A1(_04556_),
    .A2(\register_file[9][13] ),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09514_ (.A1(_04558_),
    .A2(\register_file[8][13] ),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09515_ (.A1(_04827_),
    .A2(_04828_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09516_ (.I(_04145_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09517_ (.A1(_04830_),
    .A2(\register_file[10][13] ),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09518_ (.I(_04148_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09519_ (.A1(_04832_),
    .A2(\register_file[11][13] ),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09520_ (.A1(_04831_),
    .A2(_04833_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09521_ (.A1(_04829_),
    .A2(_04834_),
    .B(_04002_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09522_ (.A1(_04630_),
    .A2(\register_file[2][13] ),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09523_ (.I(_03831_),
    .Z(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09524_ (.A1(_04837_),
    .A2(\register_file[3][13] ),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09525_ (.A1(_04633_),
    .A2(\register_file[1][13] ),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09526_ (.A1(_04836_),
    .A2(_04838_),
    .A3(_04839_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09527_ (.A1(_04840_),
    .A2(_04637_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09528_ (.A1(_04835_),
    .A2(_04841_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09529_ (.A1(_04826_),
    .A2(_04842_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09530_ (.A1(_04809_),
    .A2(_04843_),
    .B(_04641_),
    .ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09531_ (.A1(_03933_),
    .A2(\register_file[4][14] ),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09532_ (.A1(_02374_),
    .A2(_03763_),
    .B(_04844_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09533_ (.A1(_04781_),
    .A2(\register_file[6][14] ),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09534_ (.A1(_04576_),
    .A2(\register_file[7][14] ),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09535_ (.A1(_04846_),
    .A2(_04847_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09536_ (.A1(_04845_),
    .A2(_04848_),
    .B(_03962_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09537_ (.A1(_04580_),
    .A2(\register_file[25][14] ),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09538_ (.A1(_04582_),
    .A2(\register_file[24][14] ),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09539_ (.A1(_04850_),
    .A2(_04851_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09540_ (.I(_03807_),
    .Z(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09541_ (.A1(_04853_),
    .A2(\register_file[26][14] ),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09542_ (.I(_03810_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09543_ (.A1(_04855_),
    .A2(\register_file[27][14] ),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09544_ (.A1(_04854_),
    .A2(_04856_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09545_ (.A1(_04852_),
    .A2(_04857_),
    .B(_04382_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09546_ (.A1(_04849_),
    .A2(_04858_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09547_ (.A1(_04727_),
    .A2(\register_file[29][14] ),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09548_ (.A1(_04729_),
    .A2(\register_file[28][14] ),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09549_ (.A1(_04860_),
    .A2(_04861_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09550_ (.A1(_04661_),
    .A2(\register_file[30][14] ),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09551_ (.A1(_04663_),
    .A2(\register_file[31][14] ),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09552_ (.A1(_04863_),
    .A2(_04864_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09553_ (.A1(_04862_),
    .A2(_04865_),
    .B(_04183_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09554_ (.A1(_04667_),
    .A2(\register_file[13][14] ),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09555_ (.A1(_04669_),
    .A2(\register_file[12][14] ),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09556_ (.A1(_04867_),
    .A2(_04868_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09557_ (.A1(_04600_),
    .A2(\register_file[14][14] ),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09558_ (.A1(_04602_),
    .A2(\register_file[15][14] ),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09559_ (.A1(_04870_),
    .A2(_04871_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09560_ (.I(_04219_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09561_ (.A1(_04869_),
    .A2(_04872_),
    .B(_04873_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09562_ (.A1(_04866_),
    .A2(_04874_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09563_ (.A1(_04859_),
    .A2(_04875_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09564_ (.A1(_04810_),
    .A2(\register_file[9][14] ),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09565_ (.A1(_04812_),
    .A2(\register_file[8][14] ),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09566_ (.A1(_04877_),
    .A2(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09567_ (.A1(_04748_),
    .A2(\register_file[10][14] ),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09568_ (.A1(_04750_),
    .A2(\register_file[11][14] ),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09569_ (.A1(_04880_),
    .A2(_04881_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09570_ (.A1(_04879_),
    .A2(_04882_),
    .B(_04118_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09571_ (.A1(_04754_),
    .A2(\register_file[17][14] ),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(_04756_),
    .A2(\register_file[16][14] ),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09573_ (.A1(_04884_),
    .A2(_04885_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09574_ (.A1(_04689_),
    .A2(\register_file[18][14] ),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09575_ (.A1(_04691_),
    .A2(\register_file[19][14] ),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09576_ (.A1(_04887_),
    .A2(_04888_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09577_ (.A1(_04886_),
    .A2(_04889_),
    .B(_04017_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09578_ (.A1(_04883_),
    .A2(_04890_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09579_ (.I(_03897_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09580_ (.A1(_04892_),
    .A2(\register_file[21][14] ),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09581_ (.I(_03882_),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09582_ (.A1(_04894_),
    .A2(\register_file[20][14] ),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09583_ (.A1(_04893_),
    .A2(_04895_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09584_ (.A1(_04830_),
    .A2(\register_file[22][14] ),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09585_ (.A1(_04832_),
    .A2(\register_file[23][14] ),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09586_ (.A1(_04897_),
    .A2(_04898_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09587_ (.I(_03991_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09588_ (.A1(_04896_),
    .A2(_04899_),
    .B(_04900_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09589_ (.A1(_04630_),
    .A2(\register_file[2][14] ),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09590_ (.A1(_04837_),
    .A2(\register_file[3][14] ),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09591_ (.A1(_04633_),
    .A2(\register_file[1][14] ),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09592_ (.A1(_04902_),
    .A2(_04903_),
    .A3(_04904_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09593_ (.A1(_04905_),
    .A2(_04637_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09594_ (.A1(_04901_),
    .A2(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09595_ (.A1(_04891_),
    .A2(_04907_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09596_ (.A1(_04876_),
    .A2(_04908_),
    .B(_04641_),
    .ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09597_ (.A1(_04710_),
    .A2(\register_file[25][15] ),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09598_ (.A1(_04712_),
    .A2(\register_file[24][15] ),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09599_ (.A1(_04909_),
    .A2(_04910_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09600_ (.A1(_04781_),
    .A2(\register_file[26][15] ),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09601_ (.I(_03785_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09602_ (.A1(_04913_),
    .A2(\register_file[27][15] ),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09603_ (.A1(_04912_),
    .A2(_04914_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09604_ (.A1(_04911_),
    .A2(_04915_),
    .B(_03796_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09605_ (.I(_03860_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09606_ (.A1(_04917_),
    .A2(\register_file[17][15] ),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09607_ (.I(_03863_),
    .Z(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09608_ (.A1(_04919_),
    .A2(\register_file[16][15] ),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09609_ (.A1(_04918_),
    .A2(_04920_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09610_ (.A1(_04853_),
    .A2(\register_file[18][15] ),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09611_ (.A1(_04855_),
    .A2(\register_file[19][15] ),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09612_ (.A1(_04922_),
    .A2(_04923_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09613_ (.A1(_04921_),
    .A2(_04924_),
    .B(_04452_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09614_ (.A1(_04916_),
    .A2(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09615_ (.A1(_04727_),
    .A2(\register_file[13][15] ),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09616_ (.A1(_04729_),
    .A2(\register_file[12][15] ),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09617_ (.A1(_04927_),
    .A2(_04928_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09618_ (.A1(_04661_),
    .A2(\register_file[14][15] ),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09619_ (.A1(_04663_),
    .A2(\register_file[15][15] ),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09620_ (.A1(_04930_),
    .A2(_04931_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09621_ (.A1(_04929_),
    .A2(_04932_),
    .B(_03877_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09622_ (.A1(_04667_),
    .A2(\register_file[9][15] ),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09623_ (.A1(_04669_),
    .A2(\register_file[8][15] ),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09624_ (.A1(_04934_),
    .A2(_04935_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09625_ (.I(_03904_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09626_ (.A1(_04937_),
    .A2(\register_file[10][15] ),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09627_ (.I(_03907_),
    .Z(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09628_ (.A1(_04939_),
    .A2(\register_file[11][15] ),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09629_ (.A1(_04938_),
    .A2(_04940_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09630_ (.A1(_04936_),
    .A2(_04941_),
    .B(_04002_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09631_ (.A1(_04933_),
    .A2(_04942_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09632_ (.A1(_04926_),
    .A2(_04943_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09633_ (.A1(_04810_),
    .A2(\register_file[5][15] ),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09634_ (.A1(_04812_),
    .A2(\register_file[4][15] ),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09635_ (.A1(_04945_),
    .A2(_04946_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09636_ (.A1(_04748_),
    .A2(\register_file[6][15] ),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09637_ (.A1(_04750_),
    .A2(\register_file[7][15] ),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09638_ (.A1(_04948_),
    .A2(_04949_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09639_ (.A1(_04947_),
    .A2(_04950_),
    .B(_04057_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09640_ (.A1(_04754_),
    .A2(\register_file[29][15] ),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09641_ (.A1(_04756_),
    .A2(\register_file[28][15] ),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09642_ (.A1(_04952_),
    .A2(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09643_ (.A1(_04689_),
    .A2(\register_file[30][15] ),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09644_ (.A1(_04691_),
    .A2(\register_file[31][15] ),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09645_ (.A1(_04955_),
    .A2(_04956_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09646_ (.A1(_04954_),
    .A2(_04957_),
    .B(_04139_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09647_ (.A1(_04951_),
    .A2(_04958_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09648_ (.A1(_04892_),
    .A2(\register_file[21][15] ),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09649_ (.A1(_04894_),
    .A2(\register_file[20][15] ),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09650_ (.A1(_04960_),
    .A2(_04961_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09651_ (.A1(_04830_),
    .A2(\register_file[22][15] ),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09652_ (.A1(_04832_),
    .A2(\register_file[23][15] ),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09653_ (.A1(_04963_),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09654_ (.A1(_04962_),
    .A2(_04965_),
    .B(_04900_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09655_ (.I(_03916_),
    .Z(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09656_ (.A1(_04967_),
    .A2(\register_file[2][15] ),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09657_ (.A1(_04837_),
    .A2(\register_file[3][15] ),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09658_ (.I(_03776_),
    .Z(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09659_ (.A1(_04970_),
    .A2(\register_file[1][15] ),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09660_ (.A1(_04968_),
    .A2(_04969_),
    .A3(_04971_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09661_ (.I(_04636_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09662_ (.A1(_04972_),
    .A2(_04973_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09663_ (.A1(_04966_),
    .A2(_04974_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09664_ (.A1(_04959_),
    .A2(_04975_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09665_ (.I(_03934_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09666_ (.A1(_04944_),
    .A2(_04976_),
    .B(_04977_),
    .ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09667_ (.A1(_04710_),
    .A2(\register_file[25][16] ),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09668_ (.A1(_04712_),
    .A2(\register_file[24][16] ),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09669_ (.A1(_04978_),
    .A2(_04979_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09670_ (.A1(_04781_),
    .A2(\register_file[26][16] ),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09671_ (.A1(_04913_),
    .A2(\register_file[27][16] ),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09672_ (.A1(_04981_),
    .A2(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09673_ (.A1(_04980_),
    .A2(_04983_),
    .B(_03796_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09674_ (.A1(_04917_),
    .A2(\register_file[21][16] ),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09675_ (.A1(_04919_),
    .A2(\register_file[20][16] ),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09676_ (.A1(_04985_),
    .A2(_04986_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09677_ (.A1(_04853_),
    .A2(\register_file[22][16] ),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09678_ (.A1(_04855_),
    .A2(\register_file[23][16] ),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09679_ (.A1(_04988_),
    .A2(_04989_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09680_ (.A1(_04987_),
    .A2(_04990_),
    .B(_04026_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09681_ (.A1(_04984_),
    .A2(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09682_ (.A1(_04727_),
    .A2(\register_file[5][16] ),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09683_ (.A1(_04729_),
    .A2(\register_file[4][16] ),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09684_ (.A1(_04993_),
    .A2(_04994_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09685_ (.I(_04316_),
    .Z(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09686_ (.A1(_04996_),
    .A2(\register_file[6][16] ),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09687_ (.I(_04319_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09688_ (.A1(_04998_),
    .A2(\register_file[7][16] ),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09689_ (.A1(_04997_),
    .A2(_04999_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09690_ (.A1(_04995_),
    .A2(_05000_),
    .B(_04529_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09691_ (.I(_03964_),
    .Z(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09692_ (.A1(_05002_),
    .A2(\register_file[29][16] ),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09693_ (.I(_03843_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09694_ (.A1(_05004_),
    .A2(\register_file[28][16] ),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09695_ (.A1(_05003_),
    .A2(_05005_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09696_ (.A1(_04937_),
    .A2(\register_file[30][16] ),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09697_ (.A1(_04939_),
    .A2(\register_file[31][16] ),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09698_ (.A1(_05007_),
    .A2(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09699_ (.A1(_05006_),
    .A2(_05009_),
    .B(_04675_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09700_ (.A1(_05001_),
    .A2(_05010_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09701_ (.A1(_04992_),
    .A2(_05011_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09702_ (.A1(_04810_),
    .A2(\register_file[17][16] ),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09703_ (.A1(_04812_),
    .A2(\register_file[16][16] ),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09704_ (.A1(_05013_),
    .A2(_05014_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09705_ (.A1(_04748_),
    .A2(\register_file[18][16] ),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09706_ (.A1(_04750_),
    .A2(\register_file[19][16] ),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09707_ (.A1(_05016_),
    .A2(_05017_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09708_ (.A1(_05015_),
    .A2(_05018_),
    .B(_03856_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09709_ (.A1(_04754_),
    .A2(\register_file[13][16] ),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09710_ (.A1(_04756_),
    .A2(\register_file[12][16] ),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09711_ (.A1(_05020_),
    .A2(_05021_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09712_ (.I(_03886_),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09713_ (.A1(_05023_),
    .A2(\register_file[14][16] ),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09714_ (.I(_03889_),
    .Z(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09715_ (.A1(_05025_),
    .A2(\register_file[15][16] ),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09716_ (.A1(_05024_),
    .A2(_05026_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09717_ (.I(_04219_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09718_ (.A1(_05022_),
    .A2(_05027_),
    .B(_05028_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09719_ (.A1(_05019_),
    .A2(_05029_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09720_ (.A1(_04892_),
    .A2(\register_file[9][16] ),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09721_ (.A1(_04894_),
    .A2(\register_file[8][16] ),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09722_ (.A1(_05031_),
    .A2(_05032_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09723_ (.A1(_04830_),
    .A2(\register_file[10][16] ),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09724_ (.A1(_04832_),
    .A2(\register_file[11][16] ),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09725_ (.A1(_05034_),
    .A2(_05035_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09726_ (.I(_04001_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09727_ (.A1(_05033_),
    .A2(_05036_),
    .B(_05037_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09728_ (.A1(_04967_),
    .A2(\register_file[2][16] ),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09729_ (.A1(_04837_),
    .A2(\register_file[3][16] ),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09730_ (.A1(_04970_),
    .A2(\register_file[1][16] ),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09731_ (.A1(_05039_),
    .A2(_05040_),
    .A3(_05041_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09732_ (.A1(_05042_),
    .A2(_04973_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09733_ (.A1(_05038_),
    .A2(_05043_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09734_ (.A1(_05030_),
    .A2(_05044_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09735_ (.A1(_05012_),
    .A2(_05045_),
    .B(_04977_),
    .ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09736_ (.A1(_04710_),
    .A2(\register_file[9][17] ),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09737_ (.A1(_04712_),
    .A2(\register_file[8][17] ),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09738_ (.A1(_05046_),
    .A2(_05047_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09739_ (.A1(_04781_),
    .A2(\register_file[10][17] ),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09740_ (.A1(_04913_),
    .A2(\register_file[11][17] ),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09741_ (.A1(_05049_),
    .A2(_05050_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09742_ (.A1(_05048_),
    .A2(_05051_),
    .B(_04037_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09743_ (.A1(_04917_),
    .A2(\register_file[25][17] ),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09744_ (.A1(_04919_),
    .A2(\register_file[24][17] ),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09745_ (.A1(_05053_),
    .A2(_05054_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09746_ (.A1(_04853_),
    .A2(\register_file[26][17] ),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09747_ (.A1(_04855_),
    .A2(\register_file[27][17] ),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09748_ (.A1(_05056_),
    .A2(_05057_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09749_ (.A1(_05055_),
    .A2(_05058_),
    .B(_04382_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09750_ (.A1(_05052_),
    .A2(_05059_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09751_ (.I(_03820_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09752_ (.A1(_05061_),
    .A2(\register_file[17][17] ),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09753_ (.I(_03802_),
    .Z(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09754_ (.A1(_05063_),
    .A2(\register_file[16][17] ),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09755_ (.A1(_05062_),
    .A2(_05064_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09756_ (.A1(_04996_),
    .A2(\register_file[18][17] ),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09757_ (.A1(_04998_),
    .A2(\register_file[19][17] ),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09758_ (.A1(_05066_),
    .A2(_05067_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09759_ (.A1(_05065_),
    .A2(_05068_),
    .B(_04102_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09760_ (.A1(_05002_),
    .A2(\register_file[21][17] ),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09761_ (.A1(_05004_),
    .A2(\register_file[20][17] ),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09762_ (.A1(_05070_),
    .A2(_05071_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09763_ (.A1(_04937_),
    .A2(\register_file[22][17] ),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09764_ (.A1(_04939_),
    .A2(\register_file[23][17] ),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09765_ (.A1(_05073_),
    .A2(_05074_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09766_ (.A1(_05072_),
    .A2(_05075_),
    .B(_04900_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09767_ (.A1(_05069_),
    .A2(_05076_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09768_ (.A1(_05060_),
    .A2(_05077_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09769_ (.A1(_04810_),
    .A2(\register_file[5][17] ),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09770_ (.A1(_04812_),
    .A2(\register_file[4][17] ),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09771_ (.A1(_05079_),
    .A2(_05080_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09772_ (.I(_03847_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09773_ (.A1(_05082_),
    .A2(\register_file[6][17] ),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09774_ (.I(_03850_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09775_ (.A1(_05084_),
    .A2(\register_file[7][17] ),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09776_ (.A1(_05083_),
    .A2(_05085_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09777_ (.A1(_05081_),
    .A2(_05086_),
    .B(_04057_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09778_ (.I(_03765_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09779_ (.A1(_05088_),
    .A2(\register_file[29][17] ),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09780_ (.I(_04415_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09781_ (.A1(_05090_),
    .A2(\register_file[28][17] ),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09782_ (.A1(_05089_),
    .A2(_05091_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09783_ (.A1(_05023_),
    .A2(\register_file[30][17] ),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09784_ (.A1(_05025_),
    .A2(\register_file[31][17] ),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09785_ (.A1(_05093_),
    .A2(_05094_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09786_ (.A1(_05092_),
    .A2(_05095_),
    .B(_04139_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09787_ (.A1(_05087_),
    .A2(_05096_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09788_ (.A1(_04892_),
    .A2(\register_file[13][17] ),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09789_ (.A1(_04894_),
    .A2(\register_file[12][17] ),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09790_ (.A1(_05098_),
    .A2(_05099_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09791_ (.A1(_04830_),
    .A2(\register_file[14][17] ),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09792_ (.A1(_04832_),
    .A2(\register_file[15][17] ),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09793_ (.A1(_05101_),
    .A2(_05102_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09794_ (.A1(_05100_),
    .A2(_05103_),
    .B(_04220_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09795_ (.A1(_04967_),
    .A2(\register_file[2][17] ),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09796_ (.A1(_04837_),
    .A2(\register_file[3][17] ),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09797_ (.A1(_04970_),
    .A2(\register_file[1][17] ),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09798_ (.A1(_05105_),
    .A2(_05106_),
    .A3(_05107_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09799_ (.A1(_05108_),
    .A2(_04973_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09800_ (.A1(_05104_),
    .A2(_05109_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09801_ (.A1(_05097_),
    .A2(_05110_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09802_ (.A1(_05078_),
    .A2(_05111_),
    .B(_04977_),
    .ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09803_ (.I(_03766_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09804_ (.A1(_05112_),
    .A2(\register_file[21][18] ),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09805_ (.I(_03772_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09806_ (.A1(_05114_),
    .A2(\register_file[20][18] ),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09807_ (.A1(_05113_),
    .A2(_05115_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09808_ (.I(_03827_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09809_ (.A1(_05117_),
    .A2(\register_file[22][18] ),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09810_ (.A1(_04913_),
    .A2(\register_file[23][18] ),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09811_ (.A1(_05118_),
    .A2(_05119_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09812_ (.A1(_05116_),
    .A2(_05120_),
    .B(_03838_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09813_ (.A1(_04917_),
    .A2(\register_file[5][18] ),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09814_ (.A1(_04919_),
    .A2(\register_file[4][18] ),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09815_ (.A1(_05122_),
    .A2(_05123_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09816_ (.A1(_04853_),
    .A2(\register_file[6][18] ),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09817_ (.A1(_04855_),
    .A2(\register_file[7][18] ),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09818_ (.A1(_05125_),
    .A2(_05126_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09819_ (.A1(_05124_),
    .A2(_05127_),
    .B(_04655_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09820_ (.A1(_05121_),
    .A2(_05128_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09821_ (.A1(_05061_),
    .A2(\register_file[13][18] ),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09822_ (.A1(_05063_),
    .A2(\register_file[12][18] ),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09823_ (.A1(_05130_),
    .A2(_05131_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09824_ (.A1(_04996_),
    .A2(\register_file[14][18] ),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09825_ (.A1(_04998_),
    .A2(\register_file[15][18] ),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09826_ (.A1(_05133_),
    .A2(_05134_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09827_ (.A1(_05132_),
    .A2(_05135_),
    .B(_03877_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09828_ (.A1(_05002_),
    .A2(\register_file[9][18] ),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09829_ (.A1(_05004_),
    .A2(\register_file[8][18] ),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09830_ (.A1(_05137_),
    .A2(_05138_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09831_ (.A1(_04937_),
    .A2(\register_file[10][18] ),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09832_ (.A1(_04939_),
    .A2(\register_file[11][18] ),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09833_ (.A1(_05140_),
    .A2(_05141_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09834_ (.A1(_05139_),
    .A2(_05142_),
    .B(_04002_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09835_ (.A1(_05136_),
    .A2(_05143_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09836_ (.A1(_05129_),
    .A2(_05144_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09837_ (.I(_03840_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09838_ (.A1(_05146_),
    .A2(\register_file[29][18] ),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09839_ (.I(_04124_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09840_ (.A1(_05148_),
    .A2(\register_file[28][18] ),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09841_ (.A1(_05147_),
    .A2(_05149_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09842_ (.A1(_05082_),
    .A2(\register_file[30][18] ),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09843_ (.A1(_05084_),
    .A2(\register_file[31][18] ),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09844_ (.A1(_05151_),
    .A2(_05152_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09845_ (.A1(_05150_),
    .A2(_05153_),
    .B(_04675_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09846_ (.A1(_05088_),
    .A2(\register_file[17][18] ),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09847_ (.A1(_05090_),
    .A2(\register_file[16][18] ),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09848_ (.A1(_05155_),
    .A2(_05156_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09849_ (.A1(_05023_),
    .A2(\register_file[18][18] ),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09850_ (.A1(_05025_),
    .A2(\register_file[19][18] ),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09851_ (.A1(_05158_),
    .A2(_05159_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09852_ (.A1(_05157_),
    .A2(_05160_),
    .B(_04017_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09853_ (.A1(_05154_),
    .A2(_05161_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09854_ (.A1(_04892_),
    .A2(\register_file[25][18] ),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09855_ (.A1(_04894_),
    .A2(\register_file[24][18] ),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09856_ (.A1(_05163_),
    .A2(_05164_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09857_ (.I(_04145_),
    .Z(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09858_ (.A1(_05166_),
    .A2(\register_file[26][18] ),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09859_ (.I(_04148_),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09860_ (.A1(_05168_),
    .A2(\register_file[27][18] ),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09861_ (.A1(_05167_),
    .A2(_05169_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09862_ (.A1(_05165_),
    .A2(_05170_),
    .B(_04068_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09863_ (.A1(_04967_),
    .A2(\register_file[2][18] ),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09864_ (.I(_03831_),
    .Z(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09865_ (.A1(_05173_),
    .A2(\register_file[3][18] ),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09866_ (.A1(_04970_),
    .A2(\register_file[1][18] ),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09867_ (.A1(_05172_),
    .A2(_05174_),
    .A3(_05175_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09868_ (.A1(_05176_),
    .A2(_04973_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09869_ (.A1(_05171_),
    .A2(_05177_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09870_ (.A1(_05162_),
    .A2(_05178_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09871_ (.A1(_05145_),
    .A2(_05179_),
    .B(_04977_),
    .ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09872_ (.A1(_05112_),
    .A2(\register_file[13][19] ),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09873_ (.A1(_05114_),
    .A2(\register_file[12][19] ),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09874_ (.A1(_05180_),
    .A2(_05181_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09875_ (.A1(_05117_),
    .A2(\register_file[14][19] ),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09876_ (.A1(_04913_),
    .A2(\register_file[15][19] ),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09877_ (.A1(_05183_),
    .A2(_05184_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09878_ (.A1(_05182_),
    .A2(_05185_),
    .B(_04094_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09879_ (.A1(_04917_),
    .A2(\register_file[25][19] ),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09880_ (.A1(_04919_),
    .A2(\register_file[24][19] ),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09881_ (.A1(_05187_),
    .A2(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09882_ (.I(_03807_),
    .Z(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09883_ (.A1(_05190_),
    .A2(\register_file[26][19] ),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09884_ (.I(_03810_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09885_ (.A1(_05192_),
    .A2(\register_file[27][19] ),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09886_ (.A1(_05191_),
    .A2(_05193_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09887_ (.A1(_05189_),
    .A2(_05194_),
    .B(_04131_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09888_ (.A1(_05186_),
    .A2(_05195_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09889_ (.A1(_05061_),
    .A2(\register_file[5][19] ),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09890_ (.A1(_05063_),
    .A2(\register_file[4][19] ),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09891_ (.A1(_05197_),
    .A2(_05198_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09892_ (.A1(_04996_),
    .A2(\register_file[6][19] ),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09893_ (.A1(_04998_),
    .A2(\register_file[7][19] ),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09894_ (.A1(_05200_),
    .A2(_05201_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09895_ (.A1(_05199_),
    .A2(_05202_),
    .B(_04529_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09896_ (.A1(_05002_),
    .A2(\register_file[17][19] ),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09897_ (.A1(_05004_),
    .A2(\register_file[16][19] ),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09898_ (.A1(_05204_),
    .A2(_05205_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09899_ (.A1(_04937_),
    .A2(\register_file[18][19] ),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09900_ (.A1(_04939_),
    .A2(\register_file[19][19] ),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09901_ (.A1(_05207_),
    .A2(_05208_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09902_ (.A1(_05206_),
    .A2(_05209_),
    .B(_04553_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09903_ (.A1(_05203_),
    .A2(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09904_ (.A1(_05196_),
    .A2(_05211_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09905_ (.A1(_05146_),
    .A2(\register_file[29][19] ),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09906_ (.A1(_05148_),
    .A2(\register_file[28][19] ),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09907_ (.A1(_05213_),
    .A2(_05214_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09908_ (.A1(_05082_),
    .A2(\register_file[30][19] ),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09909_ (.A1(_05084_),
    .A2(\register_file[31][19] ),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09910_ (.A1(_05216_),
    .A2(_05217_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09911_ (.A1(_05215_),
    .A2(_05218_),
    .B(_04675_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09912_ (.A1(_05088_),
    .A2(\register_file[21][19] ),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09913_ (.A1(_05090_),
    .A2(\register_file[20][19] ),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09914_ (.A1(_05220_),
    .A2(_05221_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09915_ (.A1(_05023_),
    .A2(\register_file[22][19] ),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09916_ (.A1(_05025_),
    .A2(\register_file[23][19] ),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09917_ (.A1(_05223_),
    .A2(_05224_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09918_ (.A1(_05222_),
    .A2(_05225_),
    .B(_03992_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09919_ (.A1(_05219_),
    .A2(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09920_ (.I(_03879_),
    .Z(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09921_ (.A1(_05228_),
    .A2(\register_file[9][19] ),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09922_ (.I(_03882_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09923_ (.A1(_05230_),
    .A2(\register_file[8][19] ),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09924_ (.A1(_05229_),
    .A2(_05231_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09925_ (.A1(_05166_),
    .A2(\register_file[10][19] ),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09926_ (.A1(_05168_),
    .A2(\register_file[11][19] ),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09927_ (.A1(_05233_),
    .A2(_05234_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09928_ (.A1(_05232_),
    .A2(_05235_),
    .B(_05037_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09929_ (.A1(_04967_),
    .A2(\register_file[2][19] ),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09930_ (.A1(_05173_),
    .A2(\register_file[3][19] ),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09931_ (.A1(_04970_),
    .A2(\register_file[1][19] ),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09932_ (.A1(_05237_),
    .A2(_05238_),
    .A3(_05239_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09933_ (.A1(_05240_),
    .A2(_04973_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09934_ (.A1(_05236_),
    .A2(_05241_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09935_ (.A1(_05227_),
    .A2(_05242_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09936_ (.A1(_05212_),
    .A2(_05243_),
    .B(_04977_),
    .ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09937_ (.A1(_05112_),
    .A2(\register_file[29][20] ),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09938_ (.A1(_05114_),
    .A2(\register_file[28][20] ),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09939_ (.A1(_05244_),
    .A2(_05245_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09940_ (.A1(_05117_),
    .A2(\register_file[30][20] ),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09941_ (.I(_03919_),
    .Z(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09942_ (.A1(_05248_),
    .A2(\register_file[31][20] ),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09943_ (.A1(_05247_),
    .A2(_05249_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09944_ (.A1(_05246_),
    .A2(_05250_),
    .B(_03943_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09945_ (.I(_03860_),
    .Z(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09946_ (.A1(_05252_),
    .A2(\register_file[17][20] ),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09947_ (.I(_03863_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09948_ (.A1(_05254_),
    .A2(\register_file[16][20] ),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09949_ (.A1(_05253_),
    .A2(_05255_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09950_ (.A1(_05190_),
    .A2(\register_file[18][20] ),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09951_ (.A1(_05192_),
    .A2(\register_file[19][20] ),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09952_ (.A1(_05257_),
    .A2(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09953_ (.A1(_05256_),
    .A2(_05259_),
    .B(_04452_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09954_ (.A1(_05251_),
    .A2(_05260_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09955_ (.A1(_05061_),
    .A2(\register_file[9][20] ),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09956_ (.A1(_05063_),
    .A2(\register_file[8][20] ),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09957_ (.A1(_05262_),
    .A2(_05263_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09958_ (.A1(_04996_),
    .A2(\register_file[10][20] ),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09959_ (.A1(_04998_),
    .A2(\register_file[11][20] ),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09960_ (.A1(_05265_),
    .A2(_05266_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09961_ (.I(_03894_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09962_ (.A1(_05264_),
    .A2(_05267_),
    .B(_05268_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09963_ (.A1(_05002_),
    .A2(\register_file[25][20] ),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09964_ (.A1(_05004_),
    .A2(\register_file[24][20] ),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09965_ (.A1(_05270_),
    .A2(_05271_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09966_ (.I(_03904_),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09967_ (.A1(_05273_),
    .A2(\register_file[26][20] ),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09968_ (.I(_03907_),
    .Z(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09969_ (.A1(_05275_),
    .A2(\register_file[27][20] ),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09970_ (.A1(_05274_),
    .A2(_05276_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09971_ (.A1(_05272_),
    .A2(_05277_),
    .B(_04191_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09972_ (.A1(_05269_),
    .A2(_05278_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09973_ (.A1(_05261_),
    .A2(_05279_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09974_ (.A1(_05146_),
    .A2(\register_file[5][20] ),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09975_ (.A1(_05148_),
    .A2(\register_file[4][20] ),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09976_ (.A1(_05281_),
    .A2(_05282_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09977_ (.A1(_05082_),
    .A2(\register_file[6][20] ),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09978_ (.A1(_05084_),
    .A2(\register_file[7][20] ),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09979_ (.A1(_05284_),
    .A2(_05285_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09980_ (.A1(_05283_),
    .A2(_05286_),
    .B(_04057_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09981_ (.A1(_05088_),
    .A2(\register_file[13][20] ),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09982_ (.A1(_05090_),
    .A2(\register_file[12][20] ),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09983_ (.A1(_05288_),
    .A2(_05289_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09984_ (.A1(_05023_),
    .A2(\register_file[14][20] ),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09985_ (.A1(_05025_),
    .A2(\register_file[15][20] ),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09986_ (.A1(_05291_),
    .A2(_05292_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09987_ (.A1(_05290_),
    .A2(_05293_),
    .B(_05028_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09988_ (.A1(_05287_),
    .A2(_05294_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09989_ (.A1(_05228_),
    .A2(\register_file[21][20] ),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09990_ (.A1(_05230_),
    .A2(\register_file[20][20] ),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09991_ (.A1(_05296_),
    .A2(_05297_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09992_ (.A1(_05166_),
    .A2(\register_file[22][20] ),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09993_ (.A1(_05168_),
    .A2(\register_file[23][20] ),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09994_ (.A1(_05299_),
    .A2(_05300_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09995_ (.A1(_05298_),
    .A2(_05301_),
    .B(_04900_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09996_ (.I(_03779_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09997_ (.A1(_05303_),
    .A2(\register_file[2][20] ),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09998_ (.A1(_05173_),
    .A2(\register_file[3][20] ),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09999_ (.I(_03776_),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10000_ (.A1(_05306_),
    .A2(\register_file[1][20] ),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10001_ (.A1(_05304_),
    .A2(_05305_),
    .A3(_05307_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10002_ (.I(_04636_),
    .Z(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10003_ (.A1(_05308_),
    .A2(_05309_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10004_ (.A1(_05302_),
    .A2(_05310_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10005_ (.A1(_05295_),
    .A2(_05311_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10006_ (.I(_03934_),
    .Z(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10007_ (.A1(_05280_),
    .A2(_05312_),
    .B(_05313_),
    .ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10008_ (.A1(_05112_),
    .A2(\register_file[21][21] ),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10009_ (.A1(_05114_),
    .A2(\register_file[20][21] ),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10010_ (.A1(_05314_),
    .A2(_05315_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10011_ (.A1(_05117_),
    .A2(\register_file[22][21] ),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10012_ (.A1(_05248_),
    .A2(\register_file[23][21] ),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10013_ (.A1(_05317_),
    .A2(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10014_ (.A1(_05316_),
    .A2(_05319_),
    .B(_03838_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10015_ (.A1(_05252_),
    .A2(\register_file[17][21] ),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10016_ (.A1(_05254_),
    .A2(\register_file[16][21] ),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10017_ (.A1(_05321_),
    .A2(_05322_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10018_ (.A1(_05190_),
    .A2(\register_file[18][21] ),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10019_ (.A1(_05192_),
    .A2(\register_file[19][21] ),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10020_ (.A1(_05324_),
    .A2(_05325_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10021_ (.A1(_05323_),
    .A2(_05326_),
    .B(_04452_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10022_ (.A1(_05320_),
    .A2(_05327_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10023_ (.A1(_05061_),
    .A2(\register_file[5][21] ),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10024_ (.A1(_05063_),
    .A2(\register_file[4][21] ),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10025_ (.A1(_05329_),
    .A2(_05330_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10026_ (.I(_04316_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10027_ (.A1(_05332_),
    .A2(\register_file[6][21] ),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10028_ (.I(_04319_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10029_ (.A1(_05334_),
    .A2(\register_file[7][21] ),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10030_ (.A1(_05333_),
    .A2(_05335_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10031_ (.A1(_05331_),
    .A2(_05336_),
    .B(_04655_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10032_ (.I(_03964_),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10033_ (.A1(_05338_),
    .A2(\register_file[29][21] ),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10034_ (.I(_03900_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10035_ (.A1(_05340_),
    .A2(\register_file[28][21] ),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10036_ (.A1(_05339_),
    .A2(_05341_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10037_ (.A1(_05273_),
    .A2(\register_file[30][21] ),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10038_ (.A1(_05275_),
    .A2(\register_file[31][21] ),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10039_ (.A1(_05343_),
    .A2(_05344_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10040_ (.A1(_05342_),
    .A2(_05345_),
    .B(_04675_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10041_ (.A1(_05337_),
    .A2(_05346_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10042_ (.A1(_05328_),
    .A2(_05347_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10043_ (.A1(_05146_),
    .A2(\register_file[13][21] ),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10044_ (.A1(_05148_),
    .A2(\register_file[12][21] ),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10045_ (.A1(_05349_),
    .A2(_05350_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10046_ (.A1(_05082_),
    .A2(\register_file[14][21] ),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10047_ (.A1(_05084_),
    .A2(\register_file[15][21] ),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10048_ (.A1(_05352_),
    .A2(_05353_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10049_ (.A1(_05351_),
    .A2(_05354_),
    .B(_04045_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10050_ (.A1(_05088_),
    .A2(\register_file[25][21] ),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10051_ (.A1(_05090_),
    .A2(\register_file[24][21] ),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10052_ (.A1(_05356_),
    .A2(_05357_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10053_ (.I(_03778_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10054_ (.A1(_05359_),
    .A2(\register_file[26][21] ),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10055_ (.I(_03830_),
    .Z(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10056_ (.A1(_05361_),
    .A2(\register_file[27][21] ),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10057_ (.A1(_05360_),
    .A2(_05362_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10058_ (.A1(_05358_),
    .A2(_05363_),
    .B(_04486_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10059_ (.A1(_05355_),
    .A2(_05364_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10060_ (.A1(_05228_),
    .A2(\register_file[9][21] ),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10061_ (.A1(_05230_),
    .A2(\register_file[8][21] ),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10062_ (.A1(_05366_),
    .A2(_05367_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10063_ (.A1(_05166_),
    .A2(\register_file[10][21] ),
    .ZN(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10064_ (.A1(_05168_),
    .A2(\register_file[11][21] ),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10065_ (.A1(_05369_),
    .A2(_05370_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10066_ (.A1(_05368_),
    .A2(_05371_),
    .B(_05037_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10067_ (.A1(_05303_),
    .A2(\register_file[2][21] ),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10068_ (.A1(_05173_),
    .A2(\register_file[3][21] ),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10069_ (.A1(_05306_),
    .A2(\register_file[1][21] ),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10070_ (.A1(_05373_),
    .A2(_05374_),
    .A3(_05375_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10071_ (.A1(_05376_),
    .A2(_05309_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10072_ (.A1(_05372_),
    .A2(_05377_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10073_ (.A1(_05365_),
    .A2(_05378_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10074_ (.A1(_05348_),
    .A2(_05379_),
    .B(_05313_),
    .ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10075_ (.A1(_05112_),
    .A2(\register_file[17][22] ),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10076_ (.A1(_05114_),
    .A2(\register_file[16][22] ),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10077_ (.A1(_05380_),
    .A2(_05381_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10078_ (.A1(_05117_),
    .A2(\register_file[18][22] ),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10079_ (.A1(_05248_),
    .A2(\register_file[19][22] ),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10080_ (.A1(_05383_),
    .A2(_05384_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10081_ (.A1(_05382_),
    .A2(_05385_),
    .B(_04018_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10082_ (.A1(_05252_),
    .A2(\register_file[25][22] ),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10083_ (.A1(_05254_),
    .A2(\register_file[24][22] ),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10084_ (.A1(_05387_),
    .A2(_05388_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10085_ (.A1(_05190_),
    .A2(\register_file[26][22] ),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10086_ (.A1(_05192_),
    .A2(\register_file[27][22] ),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10087_ (.A1(_05390_),
    .A2(_05391_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10088_ (.A1(_05389_),
    .A2(_05392_),
    .B(_04131_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10089_ (.A1(_05386_),
    .A2(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10090_ (.I(_03799_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10091_ (.A1(_05395_),
    .A2(\register_file[29][22] ),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10092_ (.I(_03802_),
    .Z(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10093_ (.A1(_05397_),
    .A2(\register_file[28][22] ),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10094_ (.A1(_05396_),
    .A2(_05398_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10095_ (.A1(_05332_),
    .A2(\register_file[30][22] ),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10096_ (.A1(_05334_),
    .A2(\register_file[31][22] ),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10097_ (.A1(_05400_),
    .A2(_05401_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10098_ (.A1(_05399_),
    .A2(_05402_),
    .B(_04183_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10099_ (.A1(_05338_),
    .A2(\register_file[21][22] ),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10100_ (.A1(_05340_),
    .A2(\register_file[20][22] ),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10101_ (.A1(_05404_),
    .A2(_05405_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10102_ (.A1(_05273_),
    .A2(\register_file[22][22] ),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10103_ (.A1(_05275_),
    .A2(\register_file[23][22] ),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10104_ (.A1(_05407_),
    .A2(_05408_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10105_ (.A1(_05406_),
    .A2(_05409_),
    .B(_04900_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10106_ (.A1(_05403_),
    .A2(_05410_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10107_ (.A1(_05394_),
    .A2(_05411_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10108_ (.A1(_05146_),
    .A2(\register_file[5][22] ),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10109_ (.A1(_05148_),
    .A2(\register_file[4][22] ),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10110_ (.A1(_05413_),
    .A2(_05414_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10111_ (.I(_03847_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10112_ (.A1(_05416_),
    .A2(\register_file[6][22] ),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10113_ (.I(_03850_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10114_ (.A1(_05418_),
    .A2(\register_file[7][22] ),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10115_ (.A1(_05417_),
    .A2(_05419_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10116_ (.I(_03913_),
    .Z(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10117_ (.A1(_05415_),
    .A2(_05420_),
    .B(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10118_ (.I(_03765_),
    .Z(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10119_ (.A1(_05423_),
    .A2(\register_file[13][22] ),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10120_ (.I(_04415_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10121_ (.A1(_05425_),
    .A2(\register_file[12][22] ),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10122_ (.A1(_05424_),
    .A2(_05426_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10123_ (.A1(_05359_),
    .A2(\register_file[14][22] ),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10124_ (.A1(_05361_),
    .A2(\register_file[15][22] ),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10125_ (.A1(_05428_),
    .A2(_05429_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10126_ (.A1(_05427_),
    .A2(_05430_),
    .B(_03876_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10127_ (.A1(_05422_),
    .A2(_05431_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10128_ (.A1(_05228_),
    .A2(\register_file[9][22] ),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10129_ (.A1(_05230_),
    .A2(\register_file[8][22] ),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10130_ (.A1(_05433_),
    .A2(_05434_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10131_ (.A1(_05166_),
    .A2(\register_file[10][22] ),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10132_ (.A1(_05168_),
    .A2(\register_file[11][22] ),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10133_ (.A1(_05436_),
    .A2(_05437_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10134_ (.A1(_05435_),
    .A2(_05438_),
    .B(_05037_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10135_ (.A1(_05303_),
    .A2(\register_file[2][22] ),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10136_ (.A1(_05173_),
    .A2(\register_file[3][22] ),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10137_ (.A1(_05306_),
    .A2(\register_file[1][22] ),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10138_ (.A1(_05440_),
    .A2(_05441_),
    .A3(_05442_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(_05443_),
    .A2(_05309_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10140_ (.A1(_05439_),
    .A2(_05444_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10141_ (.A1(_05432_),
    .A2(_05445_),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10142_ (.A1(_05412_),
    .A2(_05446_),
    .B(_05313_),
    .ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10143_ (.I(_03766_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10144_ (.A1(_05447_),
    .A2(\register_file[29][23] ),
    .ZN(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10145_ (.I(_03823_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10146_ (.A1(_05449_),
    .A2(\register_file[28][23] ),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10147_ (.A1(_05448_),
    .A2(_05450_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10148_ (.I(_03827_),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10149_ (.A1(_05452_),
    .A2(\register_file[30][23] ),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10150_ (.A1(_05248_),
    .A2(\register_file[31][23] ),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10151_ (.A1(_05453_),
    .A2(_05454_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10152_ (.A1(_05451_),
    .A2(_05455_),
    .B(_03943_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10153_ (.A1(_05252_),
    .A2(\register_file[17][23] ),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10154_ (.A1(_05254_),
    .A2(\register_file[16][23] ),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10155_ (.A1(_05457_),
    .A2(_05458_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10156_ (.A1(_05190_),
    .A2(\register_file[18][23] ),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10157_ (.A1(_05192_),
    .A2(\register_file[19][23] ),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10158_ (.A1(_05460_),
    .A2(_05461_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10159_ (.A1(_05459_),
    .A2(_05462_),
    .B(_04452_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10160_ (.A1(_05456_),
    .A2(_05463_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10161_ (.A1(_05395_),
    .A2(\register_file[9][23] ),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10162_ (.A1(_05397_),
    .A2(\register_file[8][23] ),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10163_ (.A1(_05465_),
    .A2(_05466_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10164_ (.A1(_05332_),
    .A2(\register_file[10][23] ),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10165_ (.A1(_05334_),
    .A2(\register_file[11][23] ),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10166_ (.A1(_05468_),
    .A2(_05469_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10167_ (.A1(_05467_),
    .A2(_05470_),
    .B(_05268_),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10168_ (.A1(_05338_),
    .A2(\register_file[25][23] ),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10169_ (.A1(_05340_),
    .A2(\register_file[24][23] ),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10170_ (.A1(_05472_),
    .A2(_05473_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10171_ (.A1(_05273_),
    .A2(\register_file[26][23] ),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10172_ (.A1(_05275_),
    .A2(\register_file[27][23] ),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10173_ (.A1(_05475_),
    .A2(_05476_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10174_ (.A1(_05474_),
    .A2(_05477_),
    .B(_04191_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10175_ (.A1(_05471_),
    .A2(_05478_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10176_ (.A1(_05464_),
    .A2(_05479_),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10177_ (.I(_03840_),
    .Z(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10178_ (.A1(_05481_),
    .A2(\register_file[5][23] ),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10179_ (.I(_04124_),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10180_ (.A1(_05483_),
    .A2(\register_file[4][23] ),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10181_ (.A1(_05482_),
    .A2(_05484_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10182_ (.A1(_05416_),
    .A2(\register_file[6][23] ),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10183_ (.A1(_05418_),
    .A2(\register_file[7][23] ),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10184_ (.A1(_05486_),
    .A2(_05487_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10185_ (.A1(_05485_),
    .A2(_05488_),
    .B(_05421_),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10186_ (.A1(_05423_),
    .A2(\register_file[13][23] ),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10187_ (.A1(_05425_),
    .A2(\register_file[12][23] ),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10188_ (.A1(_05490_),
    .A2(_05491_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10189_ (.A1(_05359_),
    .A2(\register_file[14][23] ),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10190_ (.A1(_05361_),
    .A2(\register_file[15][23] ),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10191_ (.A1(_05493_),
    .A2(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10192_ (.A1(_05492_),
    .A2(_05495_),
    .B(_03876_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10193_ (.A1(_05489_),
    .A2(_05496_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10194_ (.A1(_05228_),
    .A2(\register_file[21][23] ),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10195_ (.A1(_05230_),
    .A2(\register_file[20][23] ),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10196_ (.A1(_05498_),
    .A2(_05499_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10197_ (.I(_04145_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10198_ (.A1(_05501_),
    .A2(\register_file[22][23] ),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10199_ (.I(_04148_),
    .Z(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10200_ (.A1(_05503_),
    .A2(\register_file[23][23] ),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10201_ (.A1(_05502_),
    .A2(_05504_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10202_ (.A1(_05500_),
    .A2(_05505_),
    .B(_03992_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10203_ (.A1(_05303_),
    .A2(\register_file[2][23] ),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10204_ (.I(_03831_),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10205_ (.A1(_05508_),
    .A2(\register_file[3][23] ),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10206_ (.A1(_05306_),
    .A2(\register_file[1][23] ),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10207_ (.A1(_05507_),
    .A2(_05509_),
    .A3(_05510_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10208_ (.A1(_05511_),
    .A2(_05309_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10209_ (.A1(_05506_),
    .A2(_05512_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10210_ (.A1(_05497_),
    .A2(_05513_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10211_ (.A1(_05480_),
    .A2(_05514_),
    .B(_05313_),
    .ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10212_ (.A1(_05447_),
    .A2(\register_file[17][24] ),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10213_ (.A1(_05449_),
    .A2(\register_file[16][24] ),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10214_ (.A1(_05515_),
    .A2(_05516_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10215_ (.A1(_05452_),
    .A2(\register_file[18][24] ),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10216_ (.A1(_05248_),
    .A2(\register_file[19][24] ),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10217_ (.A1(_05518_),
    .A2(_05519_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10218_ (.A1(_05517_),
    .A2(_05520_),
    .B(_04018_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10219_ (.A1(_05252_),
    .A2(\register_file[21][24] ),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10220_ (.A1(_05254_),
    .A2(\register_file[20][24] ),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10221_ (.A1(_05522_),
    .A2(_05523_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10222_ (.I(_03867_),
    .Z(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10223_ (.A1(_05525_),
    .A2(\register_file[22][24] ),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10224_ (.I(_03870_),
    .Z(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10225_ (.A1(_05527_),
    .A2(\register_file[23][24] ),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10226_ (.A1(_05526_),
    .A2(_05528_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10227_ (.A1(_05524_),
    .A2(_05529_),
    .B(_04026_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10228_ (.A1(_05521_),
    .A2(_05530_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10229_ (.A1(_05395_),
    .A2(\register_file[9][24] ),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10230_ (.A1(_05397_),
    .A2(\register_file[8][24] ),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10231_ (.A1(_05532_),
    .A2(_05533_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10232_ (.A1(_05332_),
    .A2(\register_file[10][24] ),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10233_ (.A1(_05334_),
    .A2(\register_file[11][24] ),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10234_ (.A1(_05535_),
    .A2(_05536_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10235_ (.A1(_05534_),
    .A2(_05537_),
    .B(_05268_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10236_ (.A1(_05338_),
    .A2(\register_file[13][24] ),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10237_ (.A1(_05340_),
    .A2(\register_file[12][24] ),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10238_ (.A1(_05539_),
    .A2(_05540_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10239_ (.A1(_05273_),
    .A2(\register_file[14][24] ),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10240_ (.A1(_05275_),
    .A2(\register_file[15][24] ),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10241_ (.A1(_05542_),
    .A2(_05543_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10242_ (.A1(_05541_),
    .A2(_05544_),
    .B(_04873_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10243_ (.A1(_05538_),
    .A2(_05545_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10244_ (.A1(_05531_),
    .A2(_05546_),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10245_ (.A1(_05481_),
    .A2(\register_file[5][24] ),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10246_ (.A1(_05483_),
    .A2(\register_file[4][24] ),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10247_ (.A1(_05548_),
    .A2(_05549_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10248_ (.A1(_05416_),
    .A2(\register_file[6][24] ),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10249_ (.A1(_05418_),
    .A2(\register_file[7][24] ),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10250_ (.A1(_05551_),
    .A2(_05552_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10251_ (.A1(_05550_),
    .A2(_05553_),
    .B(_05421_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10252_ (.A1(_05423_),
    .A2(\register_file[25][24] ),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10253_ (.A1(_05425_),
    .A2(\register_file[24][24] ),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10254_ (.A1(_05555_),
    .A2(_05556_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10255_ (.A1(_05359_),
    .A2(\register_file[26][24] ),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10256_ (.A1(_05361_),
    .A2(\register_file[27][24] ),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10257_ (.A1(_05558_),
    .A2(_05559_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10258_ (.A1(_05557_),
    .A2(_05560_),
    .B(_04486_),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10259_ (.A1(_05554_),
    .A2(_05561_),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10260_ (.I(_03879_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10261_ (.A1(_05563_),
    .A2(\register_file[29][24] ),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10262_ (.I(_03882_),
    .Z(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10263_ (.A1(_05565_),
    .A2(\register_file[28][24] ),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10264_ (.A1(_05564_),
    .A2(_05566_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10265_ (.A1(_05501_),
    .A2(\register_file[30][24] ),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10266_ (.A1(_05503_),
    .A2(\register_file[31][24] ),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10267_ (.A1(_05568_),
    .A2(_05569_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10268_ (.A1(_05567_),
    .A2(_05570_),
    .B(_04078_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10269_ (.A1(_05303_),
    .A2(\register_file[2][24] ),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10270_ (.A1(_05508_),
    .A2(\register_file[3][24] ),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10271_ (.A1(_05306_),
    .A2(\register_file[1][24] ),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10272_ (.A1(_05572_),
    .A2(_05573_),
    .A3(_05574_),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10273_ (.A1(_05575_),
    .A2(_05309_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10274_ (.A1(_05571_),
    .A2(_05576_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10275_ (.A1(_05562_),
    .A2(_05577_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10276_ (.A1(_05547_),
    .A2(_05578_),
    .B(_05313_),
    .ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10277_ (.A1(_05447_),
    .A2(\register_file[17][25] ),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10278_ (.A1(_05449_),
    .A2(\register_file[16][25] ),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10279_ (.A1(_05579_),
    .A2(_05580_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10280_ (.A1(_05452_),
    .A2(\register_file[18][25] ),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10281_ (.I(_03919_),
    .Z(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10282_ (.A1(_05583_),
    .A2(\register_file[19][25] ),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10283_ (.A1(_05582_),
    .A2(_05584_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10284_ (.A1(_05581_),
    .A2(_05585_),
    .B(_04018_),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10285_ (.I(_03860_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10286_ (.A1(_05587_),
    .A2(\register_file[21][25] ),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10287_ (.I(_03863_),
    .Z(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10288_ (.A1(_05589_),
    .A2(\register_file[20][25] ),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10289_ (.A1(_05588_),
    .A2(_05590_),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10290_ (.A1(_05525_),
    .A2(\register_file[22][25] ),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10291_ (.A1(_05527_),
    .A2(\register_file[23][25] ),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10292_ (.A1(_05592_),
    .A2(_05593_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10293_ (.A1(_05591_),
    .A2(_05594_),
    .B(_04026_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10294_ (.A1(_05586_),
    .A2(_05595_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10295_ (.A1(_05395_),
    .A2(\register_file[9][25] ),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10296_ (.A1(_05397_),
    .A2(\register_file[8][25] ),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10297_ (.A1(_05597_),
    .A2(_05598_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10298_ (.A1(_05332_),
    .A2(\register_file[10][25] ),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10299_ (.A1(_05334_),
    .A2(\register_file[11][25] ),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10300_ (.A1(_05600_),
    .A2(_05601_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10301_ (.A1(_05599_),
    .A2(_05602_),
    .B(_05268_),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10302_ (.A1(_05338_),
    .A2(\register_file[13][25] ),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10303_ (.A1(_05340_),
    .A2(\register_file[12][25] ),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10304_ (.A1(_05604_),
    .A2(_05605_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10305_ (.I(_03904_),
    .Z(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10306_ (.A1(_05607_),
    .A2(\register_file[14][25] ),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10307_ (.I(_03907_),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10308_ (.A1(_05609_),
    .A2(\register_file[15][25] ),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10309_ (.A1(_05608_),
    .A2(_05610_),
    .ZN(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10310_ (.A1(_05606_),
    .A2(_05611_),
    .B(_04873_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10311_ (.A1(_05603_),
    .A2(_05612_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10312_ (.A1(_05596_),
    .A2(_05613_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10313_ (.A1(_05481_),
    .A2(\register_file[5][25] ),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10314_ (.A1(_05483_),
    .A2(\register_file[4][25] ),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10315_ (.A1(_05615_),
    .A2(_05616_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10316_ (.A1(_05416_),
    .A2(\register_file[6][25] ),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10317_ (.A1(_05418_),
    .A2(\register_file[7][25] ),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10318_ (.A1(_05618_),
    .A2(_05619_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10319_ (.A1(_05617_),
    .A2(_05620_),
    .B(_05421_),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10320_ (.A1(_05423_),
    .A2(\register_file[25][25] ),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10321_ (.A1(_05425_),
    .A2(\register_file[24][25] ),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10322_ (.A1(_05622_),
    .A2(_05623_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10323_ (.A1(_05359_),
    .A2(\register_file[26][25] ),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10324_ (.A1(_05361_),
    .A2(\register_file[27][25] ),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10325_ (.A1(_05625_),
    .A2(_05626_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10326_ (.A1(_05624_),
    .A2(_05627_),
    .B(_03795_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10327_ (.A1(_05621_),
    .A2(_05628_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10328_ (.A1(_05563_),
    .A2(\register_file[29][25] ),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10329_ (.A1(_05565_),
    .A2(\register_file[28][25] ),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10330_ (.A1(_05630_),
    .A2(_05631_),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10331_ (.A1(_05501_),
    .A2(\register_file[30][25] ),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10332_ (.A1(_05503_),
    .A2(\register_file[31][25] ),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10333_ (.A1(_05633_),
    .A2(_05634_),
    .ZN(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10334_ (.A1(_05632_),
    .A2(_05635_),
    .B(_04139_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10335_ (.I(_03779_),
    .Z(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10336_ (.A1(_05637_),
    .A2(\register_file[2][25] ),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10337_ (.A1(_05508_),
    .A2(\register_file[3][25] ),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10338_ (.I(_03776_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10339_ (.A1(_05640_),
    .A2(\register_file[1][25] ),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10340_ (.A1(_05638_),
    .A2(_05639_),
    .A3(_05641_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10341_ (.I(_04636_),
    .Z(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10342_ (.A1(_05642_),
    .A2(_05643_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10343_ (.A1(_05636_),
    .A2(_05644_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10344_ (.A1(_05629_),
    .A2(_05645_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10345_ (.I(_03934_),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10346_ (.A1(_05614_),
    .A2(_05646_),
    .B(_05647_),
    .ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10347_ (.A1(_05447_),
    .A2(\register_file[17][26] ),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10348_ (.A1(_05449_),
    .A2(\register_file[16][26] ),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10349_ (.A1(_05648_),
    .A2(_05649_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10350_ (.A1(_05452_),
    .A2(\register_file[18][26] ),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10351_ (.A1(_05583_),
    .A2(\register_file[19][26] ),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10352_ (.A1(_05651_),
    .A2(_05652_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10353_ (.A1(_05650_),
    .A2(_05653_),
    .B(_04323_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10354_ (.A1(_05587_),
    .A2(\register_file[25][26] ),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10355_ (.A1(_05589_),
    .A2(\register_file[24][26] ),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10356_ (.A1(_05655_),
    .A2(_05656_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10357_ (.A1(_05525_),
    .A2(\register_file[26][26] ),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10358_ (.A1(_05527_),
    .A2(\register_file[27][26] ),
    .ZN(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10359_ (.A1(_05658_),
    .A2(_05659_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10360_ (.A1(_05657_),
    .A2(_05660_),
    .B(_04131_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10361_ (.A1(_05654_),
    .A2(_05661_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10362_ (.A1(_05395_),
    .A2(\register_file[5][26] ),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10363_ (.A1(_05397_),
    .A2(\register_file[4][26] ),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10364_ (.A1(_05663_),
    .A2(_05664_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10365_ (.I(_04316_),
    .Z(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10366_ (.A1(_05666_),
    .A2(\register_file[6][26] ),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10367_ (.I(_04319_),
    .Z(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10368_ (.A1(_05668_),
    .A2(\register_file[7][26] ),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10369_ (.A1(_05667_),
    .A2(_05669_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10370_ (.A1(_05665_),
    .A2(_05670_),
    .B(_04655_),
    .ZN(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10371_ (.I(_03897_),
    .Z(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10372_ (.A1(_05672_),
    .A2(\register_file[29][26] ),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10373_ (.I(_03900_),
    .Z(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10374_ (.A1(_05674_),
    .A2(\register_file[28][26] ),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10375_ (.A1(_05673_),
    .A2(_05675_),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10376_ (.A1(_05607_),
    .A2(\register_file[30][26] ),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10377_ (.A1(_05609_),
    .A2(\register_file[31][26] ),
    .ZN(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10378_ (.A1(_05677_),
    .A2(_05678_),
    .ZN(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10379_ (.A1(_05676_),
    .A2(_05679_),
    .B(_04078_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10380_ (.A1(_05671_),
    .A2(_05680_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10381_ (.A1(_05662_),
    .A2(_05681_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10382_ (.A1(_05481_),
    .A2(\register_file[13][26] ),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10383_ (.A1(_05483_),
    .A2(\register_file[12][26] ),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10384_ (.A1(_05683_),
    .A2(_05684_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(_05416_),
    .A2(\register_file[14][26] ),
    .ZN(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10386_ (.A1(_05418_),
    .A2(\register_file[15][26] ),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10387_ (.A1(_05686_),
    .A2(_05687_),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10388_ (.A1(_05685_),
    .A2(_05688_),
    .B(_04045_),
    .ZN(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10389_ (.A1(_05423_),
    .A2(\register_file[21][26] ),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10390_ (.A1(_05425_),
    .A2(\register_file[20][26] ),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10391_ (.A1(_05690_),
    .A2(_05691_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10392_ (.I(_03778_),
    .Z(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10393_ (.A1(_05693_),
    .A2(\register_file[22][26] ),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10394_ (.I(_03830_),
    .Z(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10395_ (.A1(_05695_),
    .A2(\register_file[23][26] ),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10396_ (.A1(_05694_),
    .A2(_05696_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10397_ (.A1(_05692_),
    .A2(_05697_),
    .B(_03992_),
    .ZN(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10398_ (.A1(_05689_),
    .A2(_05698_),
    .ZN(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10399_ (.A1(_05563_),
    .A2(\register_file[9][26] ),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10400_ (.A1(_05565_),
    .A2(\register_file[8][26] ),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10401_ (.A1(_05700_),
    .A2(_05701_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10402_ (.A1(_05501_),
    .A2(\register_file[10][26] ),
    .ZN(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10403_ (.A1(_05503_),
    .A2(\register_file[11][26] ),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10404_ (.A1(_05703_),
    .A2(_05704_),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10405_ (.A1(_05702_),
    .A2(_05705_),
    .B(_05037_),
    .ZN(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10406_ (.A1(_05637_),
    .A2(\register_file[2][26] ),
    .ZN(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10407_ (.A1(_05508_),
    .A2(\register_file[3][26] ),
    .ZN(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10408_ (.A1(_05640_),
    .A2(\register_file[1][26] ),
    .ZN(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10409_ (.A1(_05707_),
    .A2(_05708_),
    .A3(_05709_),
    .ZN(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10410_ (.A1(_05710_),
    .A2(_05643_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10411_ (.A1(_05706_),
    .A2(_05711_),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10412_ (.A1(_05699_),
    .A2(_05712_),
    .ZN(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10413_ (.A1(_05682_),
    .A2(_05713_),
    .B(_05647_),
    .ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10414_ (.A1(_05447_),
    .A2(\register_file[17][27] ),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10415_ (.A1(_05449_),
    .A2(\register_file[16][27] ),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10416_ (.A1(_05714_),
    .A2(_05715_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10417_ (.A1(_05452_),
    .A2(\register_file[18][27] ),
    .ZN(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10418_ (.A1(_05583_),
    .A2(\register_file[19][27] ),
    .ZN(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10419_ (.A1(_05717_),
    .A2(_05718_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10420_ (.A1(_05716_),
    .A2(_05719_),
    .B(_04323_),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10421_ (.A1(_05587_),
    .A2(\register_file[21][27] ),
    .ZN(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10422_ (.A1(_05589_),
    .A2(\register_file[20][27] ),
    .ZN(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10423_ (.A1(_05721_),
    .A2(_05722_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10424_ (.A1(_05525_),
    .A2(\register_file[22][27] ),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10425_ (.A1(_05527_),
    .A2(\register_file[23][27] ),
    .ZN(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10426_ (.A1(_05724_),
    .A2(_05725_),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10427_ (.A1(_05723_),
    .A2(_05726_),
    .B(_04262_),
    .ZN(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10428_ (.A1(_05720_),
    .A2(_05727_),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10429_ (.I(_03799_),
    .Z(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10430_ (.A1(_05729_),
    .A2(\register_file[9][27] ),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10431_ (.I(_03802_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10432_ (.A1(_05731_),
    .A2(\register_file[8][27] ),
    .ZN(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10433_ (.A1(_05730_),
    .A2(_05732_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10434_ (.A1(_05666_),
    .A2(\register_file[10][27] ),
    .ZN(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10435_ (.A1(_05668_),
    .A2(\register_file[11][27] ),
    .ZN(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10436_ (.A1(_05734_),
    .A2(_05735_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10437_ (.A1(_05733_),
    .A2(_05736_),
    .B(_05268_),
    .ZN(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10438_ (.A1(_05672_),
    .A2(\register_file[13][27] ),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10439_ (.A1(_05674_),
    .A2(\register_file[12][27] ),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10440_ (.A1(_05738_),
    .A2(_05739_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10441_ (.A1(_05607_),
    .A2(\register_file[14][27] ),
    .ZN(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10442_ (.A1(_05609_),
    .A2(\register_file[15][27] ),
    .ZN(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10443_ (.A1(_05741_),
    .A2(_05742_),
    .ZN(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10444_ (.A1(_05740_),
    .A2(_05743_),
    .B(_04873_),
    .ZN(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10445_ (.A1(_05737_),
    .A2(_05744_),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10446_ (.A1(_05728_),
    .A2(_05745_),
    .ZN(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10447_ (.A1(_05481_),
    .A2(\register_file[5][27] ),
    .ZN(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10448_ (.A1(_05483_),
    .A2(\register_file[4][27] ),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10449_ (.A1(_05747_),
    .A2(_05748_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10450_ (.I(_03847_),
    .Z(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10451_ (.A1(_05750_),
    .A2(\register_file[6][27] ),
    .ZN(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10452_ (.I(_03850_),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10453_ (.A1(_05752_),
    .A2(\register_file[7][27] ),
    .ZN(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10454_ (.A1(_05751_),
    .A2(_05753_),
    .ZN(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10455_ (.A1(_05749_),
    .A2(_05754_),
    .B(_05421_),
    .ZN(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10456_ (.I(_03765_),
    .Z(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10457_ (.A1(_05756_),
    .A2(\register_file[29][27] ),
    .ZN(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10458_ (.I(_04415_),
    .Z(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10459_ (.A1(_05758_),
    .A2(\register_file[28][27] ),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10460_ (.A1(_05757_),
    .A2(_05759_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10461_ (.A1(_05693_),
    .A2(\register_file[30][27] ),
    .ZN(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10462_ (.A1(_05695_),
    .A2(\register_file[31][27] ),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10463_ (.A1(_05761_),
    .A2(_05762_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10464_ (.A1(_05760_),
    .A2(_05763_),
    .B(_03816_),
    .ZN(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10465_ (.A1(_05755_),
    .A2(_05764_),
    .ZN(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10466_ (.A1(_05563_),
    .A2(\register_file[25][27] ),
    .ZN(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10467_ (.A1(_05565_),
    .A2(\register_file[24][27] ),
    .ZN(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10468_ (.A1(_05766_),
    .A2(_05767_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10469_ (.A1(_05501_),
    .A2(\register_file[26][27] ),
    .ZN(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10470_ (.A1(_05503_),
    .A2(\register_file[27][27] ),
    .ZN(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10471_ (.A1(_05769_),
    .A2(_05770_),
    .ZN(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10472_ (.A1(_05768_),
    .A2(_05771_),
    .B(_04068_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10473_ (.A1(_05637_),
    .A2(\register_file[2][27] ),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10474_ (.A1(_05508_),
    .A2(\register_file[3][27] ),
    .ZN(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10475_ (.A1(_05640_),
    .A2(\register_file[1][27] ),
    .ZN(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10476_ (.A1(_05773_),
    .A2(_05774_),
    .A3(_05775_),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10477_ (.A1(_05776_),
    .A2(_05643_),
    .ZN(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10478_ (.A1(_05772_),
    .A2(_05777_),
    .ZN(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10479_ (.A1(_05765_),
    .A2(_05778_),
    .ZN(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10480_ (.A1(_05746_),
    .A2(_05779_),
    .B(_05647_),
    .ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10481_ (.A1(_03821_),
    .A2(\register_file[17][28] ),
    .ZN(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10482_ (.A1(_03824_),
    .A2(\register_file[16][28] ),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10483_ (.A1(_05780_),
    .A2(_05781_),
    .ZN(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10484_ (.A1(_03828_),
    .A2(\register_file[18][28] ),
    .ZN(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10485_ (.A1(_05583_),
    .A2(\register_file[19][28] ),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10486_ (.A1(_05783_),
    .A2(_05784_),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10487_ (.A1(_05782_),
    .A2(_05785_),
    .B(_04323_),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10488_ (.A1(_05587_),
    .A2(\register_file[21][28] ),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10489_ (.A1(_05589_),
    .A2(\register_file[20][28] ),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10490_ (.A1(_05787_),
    .A2(_05788_),
    .ZN(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10491_ (.A1(_05525_),
    .A2(\register_file[22][28] ),
    .ZN(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10492_ (.A1(_05527_),
    .A2(\register_file[23][28] ),
    .ZN(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10493_ (.A1(_05790_),
    .A2(_05791_),
    .ZN(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10494_ (.A1(_05789_),
    .A2(_05792_),
    .B(_04262_),
    .ZN(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10495_ (.A1(_05786_),
    .A2(_05793_),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10496_ (.A1(_05729_),
    .A2(\register_file[5][28] ),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10497_ (.A1(_05731_),
    .A2(\register_file[4][28] ),
    .ZN(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10498_ (.A1(_05795_),
    .A2(_05796_),
    .ZN(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10499_ (.A1(_05666_),
    .A2(\register_file[6][28] ),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10500_ (.A1(_05668_),
    .A2(\register_file[7][28] ),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10501_ (.A1(_05798_),
    .A2(_05799_),
    .ZN(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10502_ (.A1(_05797_),
    .A2(_05800_),
    .B(_04655_),
    .ZN(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10503_ (.A1(_05672_),
    .A2(\register_file[25][28] ),
    .ZN(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10504_ (.A1(_05674_),
    .A2(\register_file[24][28] ),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10505_ (.A1(_05802_),
    .A2(_05803_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10506_ (.A1(_05607_),
    .A2(\register_file[26][28] ),
    .ZN(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10507_ (.A1(_05609_),
    .A2(\register_file[27][28] ),
    .ZN(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10508_ (.A1(_05805_),
    .A2(_05806_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10509_ (.A1(_05804_),
    .A2(_05807_),
    .B(_04191_),
    .ZN(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10510_ (.A1(_05801_),
    .A2(_05808_),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10511_ (.A1(_05794_),
    .A2(_05809_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10512_ (.A1(_03841_),
    .A2(\register_file[9][28] ),
    .ZN(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10513_ (.A1(_03844_),
    .A2(\register_file[8][28] ),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10514_ (.A1(_05811_),
    .A2(_05812_),
    .ZN(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10515_ (.A1(_05750_),
    .A2(\register_file[10][28] ),
    .ZN(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10516_ (.A1(_05752_),
    .A2(\register_file[11][28] ),
    .ZN(_05815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10517_ (.A1(_05814_),
    .A2(_05815_),
    .ZN(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10518_ (.A1(_05813_),
    .A2(_05816_),
    .B(_04118_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10519_ (.A1(_05756_),
    .A2(\register_file[29][28] ),
    .ZN(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10520_ (.A1(_05758_),
    .A2(\register_file[28][28] ),
    .ZN(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10521_ (.A1(_05818_),
    .A2(_05819_),
    .ZN(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10522_ (.A1(_05693_),
    .A2(\register_file[30][28] ),
    .ZN(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10523_ (.A1(_05695_),
    .A2(\register_file[31][28] ),
    .ZN(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10524_ (.A1(_05821_),
    .A2(_05822_),
    .ZN(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10525_ (.A1(_05820_),
    .A2(_05823_),
    .B(_03816_),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10526_ (.A1(_05817_),
    .A2(_05824_),
    .ZN(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10527_ (.A1(_05563_),
    .A2(\register_file[13][28] ),
    .ZN(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10528_ (.A1(_05565_),
    .A2(\register_file[12][28] ),
    .ZN(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10529_ (.A1(_05826_),
    .A2(_05827_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10530_ (.A1(_03887_),
    .A2(\register_file[14][28] ),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10531_ (.A1(_03890_),
    .A2(\register_file[15][28] ),
    .ZN(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10532_ (.A1(_05829_),
    .A2(_05830_),
    .ZN(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10533_ (.A1(_05828_),
    .A2(_05831_),
    .B(_05028_),
    .ZN(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10534_ (.A1(_05637_),
    .A2(\register_file[2][28] ),
    .ZN(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10535_ (.A1(_03832_),
    .A2(\register_file[3][28] ),
    .ZN(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10536_ (.A1(_05640_),
    .A2(\register_file[1][28] ),
    .ZN(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10537_ (.A1(_05833_),
    .A2(_05834_),
    .A3(_05835_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10538_ (.A1(_05836_),
    .A2(_05643_),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10539_ (.A1(_05832_),
    .A2(_05837_),
    .ZN(_05838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10540_ (.A1(_05825_),
    .A2(_05838_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10541_ (.A1(_05810_),
    .A2(_05839_),
    .B(_05647_),
    .ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10542_ (.A1(_03821_),
    .A2(\register_file[29][29] ),
    .ZN(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10543_ (.A1(_03824_),
    .A2(\register_file[28][29] ),
    .ZN(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10544_ (.A1(_05840_),
    .A2(_05841_),
    .ZN(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10545_ (.A1(_03828_),
    .A2(\register_file[30][29] ),
    .ZN(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10546_ (.A1(_05583_),
    .A2(\register_file[31][29] ),
    .ZN(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10547_ (.A1(_05843_),
    .A2(_05844_),
    .ZN(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10548_ (.A1(_05842_),
    .A2(_05845_),
    .B(_04183_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10549_ (.A1(_05587_),
    .A2(\register_file[17][29] ),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10550_ (.A1(_05589_),
    .A2(\register_file[16][29] ),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10551_ (.A1(_05847_),
    .A2(_05848_),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10552_ (.A1(_03868_),
    .A2(\register_file[18][29] ),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10553_ (.A1(_03871_),
    .A2(\register_file[19][29] ),
    .ZN(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10554_ (.A1(_05850_),
    .A2(_05851_),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10555_ (.A1(_05849_),
    .A2(_05852_),
    .B(_03856_),
    .ZN(_05853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10556_ (.A1(_05846_),
    .A2(_05853_),
    .ZN(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10557_ (.A1(_05729_),
    .A2(\register_file[9][29] ),
    .ZN(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10558_ (.A1(_05731_),
    .A2(\register_file[8][29] ),
    .ZN(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10559_ (.A1(_05855_),
    .A2(_05856_),
    .ZN(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10560_ (.A1(_05666_),
    .A2(\register_file[10][29] ),
    .ZN(_05858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10561_ (.A1(_05668_),
    .A2(\register_file[11][29] ),
    .ZN(_05859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10562_ (.A1(_05858_),
    .A2(_05859_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10563_ (.A1(_05857_),
    .A2(_05860_),
    .B(_04201_),
    .ZN(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10564_ (.A1(_05672_),
    .A2(\register_file[13][29] ),
    .ZN(_05862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10565_ (.A1(_05674_),
    .A2(\register_file[12][29] ),
    .ZN(_05863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10566_ (.A1(_05862_),
    .A2(_05863_),
    .ZN(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10567_ (.A1(_05607_),
    .A2(\register_file[14][29] ),
    .ZN(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10568_ (.A1(_05609_),
    .A2(\register_file[15][29] ),
    .ZN(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10569_ (.A1(_05865_),
    .A2(_05866_),
    .ZN(_05867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10570_ (.A1(_05864_),
    .A2(_05867_),
    .B(_04873_),
    .ZN(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10571_ (.A1(_05861_),
    .A2(_05868_),
    .ZN(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10572_ (.A1(_05854_),
    .A2(_05869_),
    .ZN(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10573_ (.A1(_03841_),
    .A2(\register_file[25][29] ),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10574_ (.A1(_03844_),
    .A2(\register_file[24][29] ),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10575_ (.A1(_05871_),
    .A2(_05872_),
    .ZN(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10576_ (.A1(_05750_),
    .A2(\register_file[26][29] ),
    .ZN(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10577_ (.A1(_05752_),
    .A2(\register_file[27][29] ),
    .ZN(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10578_ (.A1(_05874_),
    .A2(_05875_),
    .ZN(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10579_ (.A1(_05873_),
    .A2(_05876_),
    .B(_04191_),
    .ZN(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10580_ (.A1(_05756_),
    .A2(\register_file[21][29] ),
    .ZN(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10581_ (.A1(_05758_),
    .A2(\register_file[20][29] ),
    .ZN(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10582_ (.A1(_05878_),
    .A2(_05879_),
    .ZN(_05880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10583_ (.A1(_05693_),
    .A2(\register_file[22][29] ),
    .ZN(_05881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10584_ (.A1(_05695_),
    .A2(\register_file[23][29] ),
    .ZN(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10585_ (.A1(_05881_),
    .A2(_05882_),
    .ZN(_05883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10586_ (.A1(_05880_),
    .A2(_05883_),
    .B(_03837_),
    .ZN(_05884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10587_ (.A1(_05877_),
    .A2(_05884_),
    .ZN(_05885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10588_ (.A1(_03880_),
    .A2(\register_file[5][29] ),
    .ZN(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10589_ (.A1(_03883_),
    .A2(\register_file[4][29] ),
    .ZN(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10590_ (.A1(_05886_),
    .A2(_05887_),
    .ZN(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10591_ (.A1(_03887_),
    .A2(\register_file[6][29] ),
    .ZN(_05889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10592_ (.A1(_03890_),
    .A2(\register_file[7][29] ),
    .ZN(_05890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10593_ (.A1(_05889_),
    .A2(_05890_),
    .ZN(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10594_ (.A1(_05888_),
    .A2(_05891_),
    .B(_03961_),
    .ZN(_05892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10595_ (.A1(_05637_),
    .A2(\register_file[2][29] ),
    .ZN(_05893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10596_ (.A1(_03832_),
    .A2(\register_file[3][29] ),
    .ZN(_05894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10597_ (.A1(_05640_),
    .A2(\register_file[1][29] ),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10598_ (.A1(_05893_),
    .A2(_05894_),
    .A3(_05895_),
    .ZN(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10599_ (.A1(_05896_),
    .A2(_05643_),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10600_ (.A1(_05892_),
    .A2(_05897_),
    .ZN(_05898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10601_ (.A1(_05885_),
    .A2(_05898_),
    .ZN(_05899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10602_ (.A1(_05870_),
    .A2(_05899_),
    .B(_05647_),
    .ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10603_ (.A1(_03821_),
    .A2(\register_file[9][30] ),
    .ZN(_05900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10604_ (.A1(_03824_),
    .A2(\register_file[8][30] ),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10605_ (.A1(_05900_),
    .A2(_05901_),
    .ZN(_05902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10606_ (.A1(_03828_),
    .A2(\register_file[10][30] ),
    .ZN(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10607_ (.A1(_03920_),
    .A2(\register_file[11][30] ),
    .ZN(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10608_ (.A1(_05903_),
    .A2(_05904_),
    .ZN(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10609_ (.A1(_05902_),
    .A2(_05905_),
    .B(_04037_),
    .ZN(_05906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10610_ (.A1(_03861_),
    .A2(\register_file[25][30] ),
    .ZN(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10611_ (.A1(_03864_),
    .A2(\register_file[24][30] ),
    .ZN(_05908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10612_ (.A1(_05907_),
    .A2(_05908_),
    .ZN(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10613_ (.A1(_03868_),
    .A2(\register_file[26][30] ),
    .ZN(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10614_ (.A1(_03871_),
    .A2(\register_file[27][30] ),
    .ZN(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10615_ (.A1(_05910_),
    .A2(_05911_),
    .ZN(_05912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10616_ (.A1(_05909_),
    .A2(_05912_),
    .B(_04131_),
    .ZN(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10617_ (.A1(_05906_),
    .A2(_05913_),
    .ZN(_05914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10618_ (.A1(_05729_),
    .A2(\register_file[29][30] ),
    .ZN(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10619_ (.A1(_05731_),
    .A2(\register_file[28][30] ),
    .ZN(_05916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10620_ (.A1(_05915_),
    .A2(_05916_),
    .ZN(_05917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10621_ (.A1(_05666_),
    .A2(\register_file[30][30] ),
    .ZN(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10622_ (.A1(_05668_),
    .A2(\register_file[31][30] ),
    .ZN(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10623_ (.A1(_05918_),
    .A2(_05919_),
    .ZN(_05920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10624_ (.A1(_05917_),
    .A2(_05920_),
    .B(_04183_),
    .ZN(_05921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10625_ (.A1(_05672_),
    .A2(\register_file[17][30] ),
    .ZN(_05922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10626_ (.A1(_05674_),
    .A2(\register_file[16][30] ),
    .ZN(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10627_ (.A1(_05922_),
    .A2(_05923_),
    .ZN(_05924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10628_ (.A1(_03905_),
    .A2(\register_file[18][30] ),
    .ZN(_05925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10629_ (.A1(_03908_),
    .A2(\register_file[19][30] ),
    .ZN(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10630_ (.A1(_05925_),
    .A2(_05926_),
    .ZN(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10631_ (.A1(_05924_),
    .A2(_05927_),
    .B(_04553_),
    .ZN(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10632_ (.A1(_05921_),
    .A2(_05928_),
    .ZN(_05929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10633_ (.A1(_05914_),
    .A2(_05929_),
    .ZN(_05930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10634_ (.A1(_03841_),
    .A2(\register_file[5][30] ),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10635_ (.A1(_03844_),
    .A2(\register_file[4][30] ),
    .ZN(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10636_ (.A1(_05931_),
    .A2(_05932_),
    .ZN(_05933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10637_ (.A1(_05750_),
    .A2(\register_file[6][30] ),
    .ZN(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10638_ (.A1(_05752_),
    .A2(\register_file[7][30] ),
    .ZN(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10639_ (.A1(_05934_),
    .A2(_05935_),
    .ZN(_05936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10640_ (.A1(_05933_),
    .A2(_05936_),
    .B(_03914_),
    .ZN(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10641_ (.A1(_05756_),
    .A2(\register_file[21][30] ),
    .ZN(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10642_ (.A1(_05758_),
    .A2(\register_file[20][30] ),
    .ZN(_05939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10643_ (.A1(_05938_),
    .A2(_05939_),
    .ZN(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10644_ (.A1(_05693_),
    .A2(\register_file[22][30] ),
    .ZN(_05941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10645_ (.A1(_05695_),
    .A2(\register_file[23][30] ),
    .ZN(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10646_ (.A1(_05941_),
    .A2(_05942_),
    .ZN(_05943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10647_ (.A1(_05940_),
    .A2(_05943_),
    .B(_03837_),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10648_ (.A1(_05937_),
    .A2(_05944_),
    .ZN(_05945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10649_ (.A1(_03880_),
    .A2(\register_file[13][30] ),
    .ZN(_05946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10650_ (.A1(_03883_),
    .A2(\register_file[12][30] ),
    .ZN(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(_05946_),
    .A2(_05947_),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10652_ (.A1(_03887_),
    .A2(\register_file[14][30] ),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10653_ (.A1(_03890_),
    .A2(\register_file[15][30] ),
    .ZN(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10654_ (.A1(_05949_),
    .A2(_05950_),
    .ZN(_05951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10655_ (.A1(_05948_),
    .A2(_05951_),
    .B(_05028_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10656_ (.A1(_03780_),
    .A2(\register_file[2][30] ),
    .ZN(_05953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10657_ (.A1(_03832_),
    .A2(\register_file[3][30] ),
    .ZN(_05954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10658_ (.A1(_03922_),
    .A2(\register_file[1][30] ),
    .ZN(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10659_ (.A1(_05953_),
    .A2(_05954_),
    .A3(_05955_),
    .ZN(_05956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10660_ (.A1(_05956_),
    .A2(_03928_),
    .ZN(_05957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10661_ (.A1(_05952_),
    .A2(_05957_),
    .ZN(_05958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10662_ (.A1(_05945_),
    .A2(_05958_),
    .ZN(_05959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10663_ (.A1(_05930_),
    .A2(_05959_),
    .B(_03935_),
    .ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10664_ (.A1(_03933_),
    .A2(\register_file[8][31] ),
    .ZN(_05960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10665_ (.A1(_03703_),
    .A2(_03763_),
    .B(_05960_),
    .ZN(_05961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10666_ (.A1(_03828_),
    .A2(\register_file[10][31] ),
    .ZN(_05962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10667_ (.A1(_03920_),
    .A2(\register_file[11][31] ),
    .ZN(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10668_ (.A1(_05962_),
    .A2(_05963_),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10669_ (.A1(_05961_),
    .A2(_05964_),
    .B(_04037_),
    .ZN(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10670_ (.A1(_03861_),
    .A2(\register_file[21][31] ),
    .ZN(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10671_ (.A1(_03864_),
    .A2(\register_file[20][31] ),
    .ZN(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10672_ (.A1(_05966_),
    .A2(_05967_),
    .ZN(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10673_ (.A1(_03868_),
    .A2(\register_file[22][31] ),
    .ZN(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10674_ (.A1(_03871_),
    .A2(\register_file[23][31] ),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10675_ (.A1(_05969_),
    .A2(_05970_),
    .ZN(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10676_ (.A1(_05968_),
    .A2(_05971_),
    .B(_04262_),
    .ZN(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10677_ (.A1(_05965_),
    .A2(_05972_),
    .ZN(_05973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10678_ (.A1(_05729_),
    .A2(\register_file[29][31] ),
    .ZN(_05974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10679_ (.A1(_05731_),
    .A2(\register_file[28][31] ),
    .ZN(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10680_ (.A1(_05974_),
    .A2(_05975_),
    .ZN(_05976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10681_ (.A1(_03808_),
    .A2(\register_file[30][31] ),
    .ZN(_05977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10682_ (.A1(_03811_),
    .A2(\register_file[31][31] ),
    .ZN(_05978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10683_ (.A1(_05977_),
    .A2(_05978_),
    .ZN(_05979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10684_ (.A1(_05976_),
    .A2(_05979_),
    .B(_03817_),
    .ZN(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10685_ (.A1(_03898_),
    .A2(\register_file[17][31] ),
    .ZN(_05981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10686_ (.A1(_03901_),
    .A2(\register_file[16][31] ),
    .ZN(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10687_ (.A1(_05981_),
    .A2(_05982_),
    .ZN(_05983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10688_ (.A1(_03905_),
    .A2(\register_file[18][31] ),
    .ZN(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10689_ (.A1(_03908_),
    .A2(\register_file[19][31] ),
    .ZN(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10690_ (.A1(_05984_),
    .A2(_05985_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10691_ (.A1(_05983_),
    .A2(_05986_),
    .B(_04553_),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10692_ (.A1(_05980_),
    .A2(_05987_),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10693_ (.A1(_05973_),
    .A2(_05988_),
    .ZN(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10694_ (.A1(_03841_),
    .A2(\register_file[5][31] ),
    .ZN(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10695_ (.A1(_03844_),
    .A2(\register_file[4][31] ),
    .ZN(_05991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10696_ (.A1(_05990_),
    .A2(_05991_),
    .ZN(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10697_ (.A1(_05750_),
    .A2(\register_file[6][31] ),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10698_ (.A1(_05752_),
    .A2(\register_file[7][31] ),
    .ZN(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10699_ (.A1(_05993_),
    .A2(_05994_),
    .ZN(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10700_ (.A1(_05992_),
    .A2(_05995_),
    .B(_03914_),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10701_ (.A1(_05756_),
    .A2(\register_file[25][31] ),
    .ZN(_05997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10702_ (.A1(_05758_),
    .A2(\register_file[24][31] ),
    .ZN(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10703_ (.A1(_05997_),
    .A2(_05998_),
    .ZN(_05999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10704_ (.A1(_03916_),
    .A2(\register_file[26][31] ),
    .ZN(_06000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10705_ (.A1(_03785_),
    .A2(\register_file[27][31] ),
    .ZN(_06001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10706_ (.A1(_06000_),
    .A2(_06001_),
    .ZN(_06002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10707_ (.A1(_05999_),
    .A2(_06002_),
    .B(_03795_),
    .ZN(_06003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10708_ (.A1(_05996_),
    .A2(_06003_),
    .ZN(_06004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10709_ (.A1(_03880_),
    .A2(\register_file[13][31] ),
    .ZN(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10710_ (.A1(_03883_),
    .A2(\register_file[12][31] ),
    .ZN(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10711_ (.A1(_06005_),
    .A2(_06006_),
    .ZN(_06007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10712_ (.A1(_03887_),
    .A2(\register_file[14][31] ),
    .ZN(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10713_ (.A1(_03890_),
    .A2(\register_file[15][31] ),
    .ZN(_06009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10714_ (.A1(_06008_),
    .A2(_06009_),
    .ZN(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10715_ (.A1(_06007_),
    .A2(_06010_),
    .B(_05028_),
    .ZN(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10716_ (.A1(_03780_),
    .A2(\register_file[2][31] ),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10717_ (.A1(_03832_),
    .A2(\register_file[3][31] ),
    .ZN(_06013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10718_ (.A1(_03922_),
    .A2(\register_file[1][31] ),
    .ZN(_06014_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10719_ (.A1(_06012_),
    .A2(_06013_),
    .A3(_06014_),
    .ZN(_06015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10720_ (.A1(_06015_),
    .A2(_03928_),
    .ZN(_06016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10721_ (.A1(_06011_),
    .A2(_06016_),
    .ZN(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10722_ (.A1(_06004_),
    .A2(_06017_),
    .ZN(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10723_ (.A1(_05989_),
    .A2(_06018_),
    .B(_03935_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10724_ (.I(net11),
    .ZN(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10725_ (.I(_06019_),
    .Z(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10726_ (.I(_06020_),
    .Z(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10727_ (.A1(_03777_),
    .A2(net43),
    .ZN(_06022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10728_ (.I(_06022_),
    .ZN(_06023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10729_ (.I(_06023_),
    .Z(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10730_ (.A1(_06024_),
    .A2(_04077_),
    .ZN(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10731_ (.I(_06025_),
    .Z(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10732_ (.I(_06026_),
    .Z(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10733_ (.I(_06025_),
    .Z(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10734_ (.I(_06028_),
    .Z(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(_06029_),
    .A2(\register_file[30][0] ),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10736_ (.A1(_06021_),
    .A2(_06027_),
    .B(_06030_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10737_ (.I(net22),
    .ZN(_06031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10738_ (.I(_06031_),
    .Z(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10739_ (.I(_06032_),
    .Z(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10740_ (.A1(_06029_),
    .A2(\register_file[30][1] ),
    .ZN(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10741_ (.A1(_06033_),
    .A2(_06027_),
    .B(_06034_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10742_ (.I(net33),
    .ZN(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10743_ (.I(_06035_),
    .Z(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10744_ (.I(_06036_),
    .Z(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10745_ (.A1(_06029_),
    .A2(\register_file[30][2] ),
    .ZN(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10746_ (.A1(_06037_),
    .A2(_06027_),
    .B(_06038_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10747_ (.I(net36),
    .ZN(_06039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10748_ (.I(_06039_),
    .Z(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10749_ (.I(_06040_),
    .Z(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10750_ (.I(_06028_),
    .Z(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10751_ (.A1(_06042_),
    .A2(\register_file[30][3] ),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10752_ (.A1(_06041_),
    .A2(_06027_),
    .B(_06043_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10753_ (.I(net37),
    .ZN(_06044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10754_ (.I(_06044_),
    .Z(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10755_ (.I(_06045_),
    .Z(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10756_ (.A1(_06042_),
    .A2(\register_file[30][4] ),
    .ZN(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10757_ (.A1(_06046_),
    .A2(_06027_),
    .B(_06047_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10758_ (.I(net38),
    .ZN(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10759_ (.I(_06048_),
    .Z(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10760_ (.I(_06049_),
    .Z(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10761_ (.I(_06028_),
    .Z(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10762_ (.I(_06051_),
    .Z(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10763_ (.A1(_06042_),
    .A2(\register_file[30][5] ),
    .ZN(_06053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10764_ (.A1(_06050_),
    .A2(_06052_),
    .B(_06053_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10765_ (.I(net39),
    .ZN(_06054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10766_ (.I(_06054_),
    .Z(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10767_ (.I(_06055_),
    .Z(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10768_ (.A1(_06042_),
    .A2(\register_file[30][6] ),
    .ZN(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10769_ (.A1(_06056_),
    .A2(_06052_),
    .B(_06057_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10770_ (.I(net40),
    .ZN(_06058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10771_ (.I(_06058_),
    .Z(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10772_ (.I(_06059_),
    .Z(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(_06042_),
    .A2(\register_file[30][7] ),
    .ZN(_06061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10774_ (.A1(_06060_),
    .A2(_06052_),
    .B(_06061_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10775_ (.I(net41),
    .ZN(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10776_ (.I(_06062_),
    .Z(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10777_ (.I(_06063_),
    .Z(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10778_ (.I(_06028_),
    .Z(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(_06065_),
    .A2(\register_file[30][8] ),
    .ZN(_06066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10780_ (.A1(_06064_),
    .A2(_06052_),
    .B(_06066_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10781_ (.I(net42),
    .ZN(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10782_ (.I(_06067_),
    .Z(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10783_ (.I(_06068_),
    .Z(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10784_ (.A1(_06065_),
    .A2(\register_file[30][9] ),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10785_ (.A1(_06069_),
    .A2(_06052_),
    .B(_06070_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10786_ (.I(net12),
    .ZN(_06071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10787_ (.I(_06071_),
    .Z(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10788_ (.I(_06072_),
    .Z(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10789_ (.I(_06051_),
    .Z(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10790_ (.A1(_06065_),
    .A2(\register_file[30][10] ),
    .ZN(_06075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10791_ (.A1(_06073_),
    .A2(_06074_),
    .B(_06075_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10792_ (.I(net13),
    .ZN(_06076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10793_ (.I(_06076_),
    .Z(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10794_ (.I(_06077_),
    .Z(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10795_ (.A1(_06065_),
    .A2(\register_file[30][11] ),
    .ZN(_06079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10796_ (.A1(_06078_),
    .A2(_06074_),
    .B(_06079_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10797_ (.I(net14),
    .ZN(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10798_ (.I(_06080_),
    .Z(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10799_ (.I(_06081_),
    .Z(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10800_ (.A1(_06065_),
    .A2(\register_file[30][12] ),
    .ZN(_06083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10801_ (.A1(_06082_),
    .A2(_06074_),
    .B(_06083_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10802_ (.I(net15),
    .ZN(_06084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10803_ (.I(_06084_),
    .Z(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10804_ (.I(_06085_),
    .Z(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10805_ (.I(_06028_),
    .Z(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10806_ (.A1(_06087_),
    .A2(\register_file[30][13] ),
    .ZN(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10807_ (.A1(_06086_),
    .A2(_06074_),
    .B(_06088_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10808_ (.I(net16),
    .ZN(_06089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10809_ (.I(_06089_),
    .Z(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10810_ (.I(_06090_),
    .Z(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10811_ (.A1(_06087_),
    .A2(\register_file[30][14] ),
    .ZN(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10812_ (.A1(_06091_),
    .A2(_06074_),
    .B(_06092_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10813_ (.I(net17),
    .ZN(_06093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10814_ (.I(_06093_),
    .Z(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10815_ (.I(_06094_),
    .Z(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10816_ (.I(_06051_),
    .Z(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10817_ (.A1(_06087_),
    .A2(\register_file[30][15] ),
    .ZN(_06097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10818_ (.A1(_06095_),
    .A2(_06096_),
    .B(_06097_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10819_ (.I(net18),
    .ZN(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10820_ (.I(_06098_),
    .Z(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10821_ (.I(_06099_),
    .Z(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10822_ (.A1(_06087_),
    .A2(\register_file[30][16] ),
    .ZN(_06101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10823_ (.A1(_06100_),
    .A2(_06096_),
    .B(_06101_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10824_ (.I(net19),
    .ZN(_06102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10825_ (.I(_06102_),
    .Z(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10826_ (.I(_06103_),
    .Z(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10827_ (.A1(_06087_),
    .A2(\register_file[30][17] ),
    .ZN(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10828_ (.A1(_06104_),
    .A2(_06096_),
    .B(_06105_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10829_ (.I(net20),
    .ZN(_06106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10830_ (.I(_06106_),
    .Z(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10831_ (.I(_06107_),
    .Z(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10832_ (.I(_06025_),
    .Z(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10833_ (.A1(_06109_),
    .A2(\register_file[30][18] ),
    .ZN(_06110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10834_ (.A1(_06108_),
    .A2(_06096_),
    .B(_06110_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10835_ (.I(net21),
    .ZN(_06111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10836_ (.I(_06111_),
    .Z(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10837_ (.I(_06112_),
    .Z(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10838_ (.A1(_06109_),
    .A2(\register_file[30][19] ),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10839_ (.A1(_06113_),
    .A2(_06096_),
    .B(_06114_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10840_ (.I(net23),
    .ZN(_06115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10841_ (.I(_06115_),
    .Z(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10842_ (.I(_06116_),
    .Z(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10843_ (.I(_06051_),
    .Z(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10844_ (.A1(_06109_),
    .A2(\register_file[30][20] ),
    .ZN(_06119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10845_ (.A1(_06117_),
    .A2(_06118_),
    .B(_06119_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10846_ (.I(net24),
    .ZN(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10847_ (.I(_06120_),
    .Z(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10848_ (.I(_06121_),
    .Z(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10849_ (.A1(_06109_),
    .A2(\register_file[30][21] ),
    .ZN(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10850_ (.A1(_06122_),
    .A2(_06118_),
    .B(_06123_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10851_ (.I(net25),
    .ZN(_06124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10852_ (.I(_06124_),
    .Z(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10853_ (.I(_06125_),
    .Z(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10854_ (.A1(_06109_),
    .A2(\register_file[30][22] ),
    .ZN(_06127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10855_ (.A1(_06126_),
    .A2(_06118_),
    .B(_06127_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10856_ (.I(net26),
    .ZN(_06128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10857_ (.I(_06128_),
    .Z(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10858_ (.I(_06129_),
    .Z(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10859_ (.I(_06025_),
    .Z(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10860_ (.A1(_06131_),
    .A2(\register_file[30][23] ),
    .ZN(_06132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10861_ (.A1(_06130_),
    .A2(_06118_),
    .B(_06132_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10862_ (.I(net27),
    .ZN(_06133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10863_ (.I(_06133_),
    .Z(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10864_ (.I(_06134_),
    .Z(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10865_ (.A1(_06131_),
    .A2(\register_file[30][24] ),
    .ZN(_06136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10866_ (.A1(_06135_),
    .A2(_06118_),
    .B(_06136_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10867_ (.I(net28),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10868_ (.I(_06137_),
    .Z(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10869_ (.I(_06138_),
    .Z(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10870_ (.I(_06051_),
    .Z(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10871_ (.A1(_06131_),
    .A2(\register_file[30][25] ),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10872_ (.A1(_06139_),
    .A2(_06140_),
    .B(_06141_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10873_ (.I(net29),
    .ZN(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10874_ (.I(_06142_),
    .Z(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10875_ (.I(_06143_),
    .Z(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_06131_),
    .A2(\register_file[30][26] ),
    .ZN(_06145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10877_ (.A1(_06144_),
    .A2(_06140_),
    .B(_06145_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10878_ (.I(net30),
    .ZN(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10879_ (.I(_06146_),
    .Z(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10880_ (.I(_06147_),
    .Z(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10881_ (.A1(_06131_),
    .A2(\register_file[30][27] ),
    .ZN(_06149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10882_ (.A1(_06148_),
    .A2(_06140_),
    .B(_06149_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10883_ (.I(net31),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10884_ (.I(_06150_),
    .Z(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10885_ (.I(_06151_),
    .Z(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10886_ (.A1(_06026_),
    .A2(\register_file[30][28] ),
    .ZN(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10887_ (.A1(_06152_),
    .A2(_06140_),
    .B(_06153_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10888_ (.I(net32),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10889_ (.I(_06154_),
    .Z(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10890_ (.I(_06155_),
    .Z(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10891_ (.A1(_06026_),
    .A2(\register_file[30][29] ),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10892_ (.A1(_06156_),
    .A2(_06140_),
    .B(_06157_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10893_ (.I(net34),
    .ZN(_06158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10894_ (.I(_06158_),
    .Z(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10895_ (.I(_06159_),
    .Z(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10896_ (.A1(_06026_),
    .A2(\register_file[30][30] ),
    .ZN(_06161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10897_ (.A1(_06160_),
    .A2(_06029_),
    .B(_06161_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10898_ (.I(net35),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10899_ (.I(_06162_),
    .Z(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10900_ (.I(_06163_),
    .Z(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10901_ (.A1(_06026_),
    .A2(\register_file[30][31] ),
    .ZN(_06165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10902_ (.A1(_06164_),
    .A2(_06029_),
    .B(_06165_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10903_ (.A1(_06024_),
    .A2(_04636_),
    .ZN(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10904_ (.I(_06166_),
    .Z(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10905_ (.I(_06167_),
    .Z(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10906_ (.I(_06166_),
    .Z(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10907_ (.I(_06169_),
    .Z(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10908_ (.A1(_06170_),
    .A2(\register_file[2][0] ),
    .ZN(_06171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10909_ (.A1(_06021_),
    .A2(_06168_),
    .B(_06171_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10910_ (.A1(_06170_),
    .A2(\register_file[2][1] ),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10911_ (.A1(_06033_),
    .A2(_06168_),
    .B(_06172_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10912_ (.A1(_06170_),
    .A2(\register_file[2][2] ),
    .ZN(_06173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10913_ (.A1(_06037_),
    .A2(_06168_),
    .B(_06173_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10914_ (.I(_06169_),
    .Z(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10915_ (.A1(_06174_),
    .A2(\register_file[2][3] ),
    .ZN(_06175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10916_ (.A1(_06041_),
    .A2(_06168_),
    .B(_06175_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10917_ (.A1(_06174_),
    .A2(\register_file[2][4] ),
    .ZN(_06176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10918_ (.A1(_06046_),
    .A2(_06168_),
    .B(_06176_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10919_ (.I(_06169_),
    .Z(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10920_ (.I(_06177_),
    .Z(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10921_ (.A1(_06174_),
    .A2(\register_file[2][5] ),
    .ZN(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10922_ (.A1(_06050_),
    .A2(_06178_),
    .B(_06179_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10923_ (.A1(_06174_),
    .A2(\register_file[2][6] ),
    .ZN(_06180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10924_ (.A1(_06056_),
    .A2(_06178_),
    .B(_06180_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10925_ (.A1(_06174_),
    .A2(\register_file[2][7] ),
    .ZN(_06181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10926_ (.A1(_06060_),
    .A2(_06178_),
    .B(_06181_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10927_ (.I(_06169_),
    .Z(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10928_ (.A1(_06182_),
    .A2(\register_file[2][8] ),
    .ZN(_06183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10929_ (.A1(_06064_),
    .A2(_06178_),
    .B(_06183_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10930_ (.A1(_06182_),
    .A2(\register_file[2][9] ),
    .ZN(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10931_ (.A1(_06069_),
    .A2(_06178_),
    .B(_06184_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10932_ (.I(_06177_),
    .Z(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10933_ (.A1(_06182_),
    .A2(\register_file[2][10] ),
    .ZN(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10934_ (.A1(_06073_),
    .A2(_06185_),
    .B(_06186_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10935_ (.A1(_06182_),
    .A2(\register_file[2][11] ),
    .ZN(_06187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10936_ (.A1(_06078_),
    .A2(_06185_),
    .B(_06187_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10937_ (.A1(_06182_),
    .A2(\register_file[2][12] ),
    .ZN(_06188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10938_ (.A1(_06082_),
    .A2(_06185_),
    .B(_06188_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10939_ (.I(_06169_),
    .Z(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10940_ (.A1(_06189_),
    .A2(\register_file[2][13] ),
    .ZN(_06190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10941_ (.A1(_06086_),
    .A2(_06185_),
    .B(_06190_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10942_ (.A1(_06189_),
    .A2(\register_file[2][14] ),
    .ZN(_06191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10943_ (.A1(_06091_),
    .A2(_06185_),
    .B(_06191_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10944_ (.I(_06177_),
    .Z(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10945_ (.A1(_06189_),
    .A2(\register_file[2][15] ),
    .ZN(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10946_ (.A1(_06095_),
    .A2(_06192_),
    .B(_06193_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10947_ (.A1(_06189_),
    .A2(\register_file[2][16] ),
    .ZN(_06194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10948_ (.A1(_06100_),
    .A2(_06192_),
    .B(_06194_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10949_ (.A1(_06189_),
    .A2(\register_file[2][17] ),
    .ZN(_06195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10950_ (.A1(_06104_),
    .A2(_06192_),
    .B(_06195_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10951_ (.I(_06166_),
    .Z(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10952_ (.A1(_06196_),
    .A2(\register_file[2][18] ),
    .ZN(_06197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10953_ (.A1(_06108_),
    .A2(_06192_),
    .B(_06197_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10954_ (.A1(_06196_),
    .A2(\register_file[2][19] ),
    .ZN(_06198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10955_ (.A1(_06113_),
    .A2(_06192_),
    .B(_06198_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10956_ (.I(_06177_),
    .Z(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10957_ (.A1(_06196_),
    .A2(\register_file[2][20] ),
    .ZN(_06200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10958_ (.A1(_06117_),
    .A2(_06199_),
    .B(_06200_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10959_ (.A1(_06196_),
    .A2(\register_file[2][21] ),
    .ZN(_06201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10960_ (.A1(_06122_),
    .A2(_06199_),
    .B(_06201_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10961_ (.A1(_06196_),
    .A2(\register_file[2][22] ),
    .ZN(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10962_ (.A1(_06126_),
    .A2(_06199_),
    .B(_06202_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10963_ (.I(_06166_),
    .Z(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10964_ (.A1(_06203_),
    .A2(\register_file[2][23] ),
    .ZN(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10965_ (.A1(_06130_),
    .A2(_06199_),
    .B(_06204_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10966_ (.A1(_06203_),
    .A2(\register_file[2][24] ),
    .ZN(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10967_ (.A1(_06135_),
    .A2(_06199_),
    .B(_06205_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10968_ (.I(_06177_),
    .Z(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10969_ (.A1(_06203_),
    .A2(\register_file[2][25] ),
    .ZN(_06207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10970_ (.A1(_06139_),
    .A2(_06206_),
    .B(_06207_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10971_ (.A1(_06203_),
    .A2(\register_file[2][26] ),
    .ZN(_06208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10972_ (.A1(_06144_),
    .A2(_06206_),
    .B(_06208_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10973_ (.A1(_06203_),
    .A2(\register_file[2][27] ),
    .ZN(_06209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10974_ (.A1(_06148_),
    .A2(_06206_),
    .B(_06209_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10975_ (.A1(_06167_),
    .A2(\register_file[2][28] ),
    .ZN(_06210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10976_ (.A1(_06152_),
    .A2(_06206_),
    .B(_06210_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10977_ (.A1(_06167_),
    .A2(\register_file[2][29] ),
    .ZN(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10978_ (.A1(_06156_),
    .A2(_06206_),
    .B(_06211_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10979_ (.A1(_06167_),
    .A2(\register_file[2][30] ),
    .ZN(_06212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10980_ (.A1(_06160_),
    .A2(_06170_),
    .B(_06212_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10981_ (.A1(_06167_),
    .A2(\register_file[2][31] ),
    .ZN(_06213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10982_ (.A1(_06164_),
    .A2(_06170_),
    .B(_06213_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10983_ (.A1(_03769_),
    .A2(net43),
    .ZN(_06214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10984_ (.I(_06214_),
    .ZN(_06215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10985_ (.I(_06215_),
    .Z(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10986_ (.A1(_04077_),
    .A2(_06216_),
    .ZN(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10987_ (.I(_06217_),
    .Z(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10988_ (.I(_06218_),
    .Z(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10989_ (.I(_06217_),
    .Z(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10990_ (.I(_06220_),
    .Z(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10991_ (.A1(_06221_),
    .A2(\register_file[28][0] ),
    .ZN(_06222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10992_ (.A1(_06021_),
    .A2(_06219_),
    .B(_06222_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10993_ (.A1(_06221_),
    .A2(\register_file[28][1] ),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10994_ (.A1(_06033_),
    .A2(_06219_),
    .B(_06223_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10995_ (.A1(_06221_),
    .A2(\register_file[28][2] ),
    .ZN(_06224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10996_ (.A1(_06037_),
    .A2(_06219_),
    .B(_06224_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10997_ (.I(_06220_),
    .Z(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10998_ (.A1(_06225_),
    .A2(\register_file[28][3] ),
    .ZN(_06226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10999_ (.A1(_06041_),
    .A2(_06219_),
    .B(_06226_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11000_ (.A1(_06225_),
    .A2(\register_file[28][4] ),
    .ZN(_06227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11001_ (.A1(_06046_),
    .A2(_06219_),
    .B(_06227_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11002_ (.I(_06220_),
    .Z(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11003_ (.I(_06228_),
    .Z(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11004_ (.A1(_06225_),
    .A2(\register_file[28][5] ),
    .ZN(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11005_ (.A1(_06050_),
    .A2(_06229_),
    .B(_06230_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11006_ (.A1(_06225_),
    .A2(\register_file[28][6] ),
    .ZN(_06231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11007_ (.A1(_06056_),
    .A2(_06229_),
    .B(_06231_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11008_ (.A1(_06225_),
    .A2(\register_file[28][7] ),
    .ZN(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11009_ (.A1(_06060_),
    .A2(_06229_),
    .B(_06232_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11010_ (.I(_06220_),
    .Z(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11011_ (.A1(_06233_),
    .A2(\register_file[28][8] ),
    .ZN(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11012_ (.A1(_06064_),
    .A2(_06229_),
    .B(_06234_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11013_ (.A1(_06233_),
    .A2(\register_file[28][9] ),
    .ZN(_06235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11014_ (.A1(_06069_),
    .A2(_06229_),
    .B(_06235_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11015_ (.I(_06228_),
    .Z(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11016_ (.A1(_06233_),
    .A2(\register_file[28][10] ),
    .ZN(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11017_ (.A1(_06073_),
    .A2(_06236_),
    .B(_06237_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11018_ (.A1(_06233_),
    .A2(\register_file[28][11] ),
    .ZN(_06238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11019_ (.A1(_06078_),
    .A2(_06236_),
    .B(_06238_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11020_ (.A1(_06233_),
    .A2(\register_file[28][12] ),
    .ZN(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11021_ (.A1(_06082_),
    .A2(_06236_),
    .B(_06239_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11022_ (.I(_06220_),
    .Z(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11023_ (.A1(_06240_),
    .A2(\register_file[28][13] ),
    .ZN(_06241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11024_ (.A1(_06086_),
    .A2(_06236_),
    .B(_06241_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11025_ (.A1(_06240_),
    .A2(\register_file[28][14] ),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11026_ (.A1(_06091_),
    .A2(_06236_),
    .B(_06242_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11027_ (.I(_06228_),
    .Z(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11028_ (.A1(_06240_),
    .A2(\register_file[28][15] ),
    .ZN(_06244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11029_ (.A1(_06095_),
    .A2(_06243_),
    .B(_06244_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11030_ (.A1(_06240_),
    .A2(\register_file[28][16] ),
    .ZN(_06245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11031_ (.A1(_06100_),
    .A2(_06243_),
    .B(_06245_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11032_ (.A1(_06240_),
    .A2(\register_file[28][17] ),
    .ZN(_06246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11033_ (.A1(_06104_),
    .A2(_06243_),
    .B(_06246_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11034_ (.I(_06217_),
    .Z(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11035_ (.A1(_06247_),
    .A2(\register_file[28][18] ),
    .ZN(_06248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11036_ (.A1(_06108_),
    .A2(_06243_),
    .B(_06248_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11037_ (.A1(_06247_),
    .A2(\register_file[28][19] ),
    .ZN(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11038_ (.A1(_06113_),
    .A2(_06243_),
    .B(_06249_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11039_ (.I(_06228_),
    .Z(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11040_ (.A1(_06247_),
    .A2(\register_file[28][20] ),
    .ZN(_06251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11041_ (.A1(_06117_),
    .A2(_06250_),
    .B(_06251_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11042_ (.A1(_06247_),
    .A2(\register_file[28][21] ),
    .ZN(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11043_ (.A1(_06122_),
    .A2(_06250_),
    .B(_06252_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11044_ (.A1(_06247_),
    .A2(\register_file[28][22] ),
    .ZN(_06253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11045_ (.A1(_06126_),
    .A2(_06250_),
    .B(_06253_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11046_ (.I(_06217_),
    .Z(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11047_ (.A1(_06254_),
    .A2(\register_file[28][23] ),
    .ZN(_06255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11048_ (.A1(_06130_),
    .A2(_06250_),
    .B(_06255_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11049_ (.A1(_06254_),
    .A2(\register_file[28][24] ),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11050_ (.A1(_06135_),
    .A2(_06250_),
    .B(_06256_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11051_ (.I(_06228_),
    .Z(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11052_ (.A1(_06254_),
    .A2(\register_file[28][25] ),
    .ZN(_06258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11053_ (.A1(_06139_),
    .A2(_06257_),
    .B(_06258_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11054_ (.A1(_06254_),
    .A2(\register_file[28][26] ),
    .ZN(_06259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11055_ (.A1(_06144_),
    .A2(_06257_),
    .B(_06259_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11056_ (.A1(_06254_),
    .A2(\register_file[28][27] ),
    .ZN(_06260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11057_ (.A1(_06148_),
    .A2(_06257_),
    .B(_06260_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11058_ (.A1(_06218_),
    .A2(\register_file[28][28] ),
    .ZN(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11059_ (.A1(_06152_),
    .A2(_06257_),
    .B(_06261_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11060_ (.A1(_06218_),
    .A2(\register_file[28][29] ),
    .ZN(_06262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11061_ (.A1(_06156_),
    .A2(_06257_),
    .B(_06262_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11062_ (.A1(_06218_),
    .A2(\register_file[28][30] ),
    .ZN(_06263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11063_ (.A1(_06160_),
    .A2(_06221_),
    .B(_06263_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11064_ (.A1(_06218_),
    .A2(\register_file[28][31] ),
    .ZN(_06264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11065_ (.A1(_06164_),
    .A2(_06221_),
    .B(_06264_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11066_ (.A1(_03783_),
    .A2(net43),
    .Z(_06265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11067_ (.I(_06265_),
    .Z(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11068_ (.A1(_06266_),
    .A2(_04067_),
    .ZN(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11069_ (.I(_06267_),
    .Z(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11070_ (.I(_06268_),
    .Z(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11071_ (.I(_06267_),
    .Z(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11072_ (.I(_06270_),
    .Z(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11073_ (.A1(_06271_),
    .A2(\register_file[27][0] ),
    .ZN(_06272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11074_ (.A1(_06021_),
    .A2(_06269_),
    .B(_06272_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11075_ (.A1(_06271_),
    .A2(\register_file[27][1] ),
    .ZN(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11076_ (.A1(_06033_),
    .A2(_06269_),
    .B(_06273_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11077_ (.A1(_06271_),
    .A2(\register_file[27][2] ),
    .ZN(_06274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11078_ (.A1(_06037_),
    .A2(_06269_),
    .B(_06274_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11079_ (.I(_06270_),
    .Z(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11080_ (.A1(_06275_),
    .A2(\register_file[27][3] ),
    .ZN(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11081_ (.A1(_06041_),
    .A2(_06269_),
    .B(_06276_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11082_ (.A1(_06275_),
    .A2(\register_file[27][4] ),
    .ZN(_06277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11083_ (.A1(_06046_),
    .A2(_06269_),
    .B(_06277_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11084_ (.I(_06270_),
    .Z(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11085_ (.I(_06278_),
    .Z(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11086_ (.A1(_06275_),
    .A2(\register_file[27][5] ),
    .ZN(_06280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11087_ (.A1(_06050_),
    .A2(_06279_),
    .B(_06280_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11088_ (.A1(_06275_),
    .A2(\register_file[27][6] ),
    .ZN(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11089_ (.A1(_06056_),
    .A2(_06279_),
    .B(_06281_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11090_ (.A1(_06275_),
    .A2(\register_file[27][7] ),
    .ZN(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11091_ (.A1(_06060_),
    .A2(_06279_),
    .B(_06282_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11092_ (.I(_06270_),
    .Z(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11093_ (.A1(_06283_),
    .A2(\register_file[27][8] ),
    .ZN(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11094_ (.A1(_06064_),
    .A2(_06279_),
    .B(_06284_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11095_ (.A1(_06283_),
    .A2(\register_file[27][9] ),
    .ZN(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11096_ (.A1(_06069_),
    .A2(_06279_),
    .B(_06285_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11097_ (.I(_06278_),
    .Z(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11098_ (.A1(_06283_),
    .A2(\register_file[27][10] ),
    .ZN(_06287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11099_ (.A1(_06073_),
    .A2(_06286_),
    .B(_06287_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11100_ (.A1(_06283_),
    .A2(\register_file[27][11] ),
    .ZN(_06288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11101_ (.A1(_06078_),
    .A2(_06286_),
    .B(_06288_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11102_ (.A1(_06283_),
    .A2(\register_file[27][12] ),
    .ZN(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11103_ (.A1(_06082_),
    .A2(_06286_),
    .B(_06289_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11104_ (.I(_06270_),
    .Z(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11105_ (.A1(_06290_),
    .A2(\register_file[27][13] ),
    .ZN(_06291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11106_ (.A1(_06086_),
    .A2(_06286_),
    .B(_06291_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11107_ (.A1(_06290_),
    .A2(\register_file[27][14] ),
    .ZN(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11108_ (.A1(_06091_),
    .A2(_06286_),
    .B(_06292_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11109_ (.I(_06278_),
    .Z(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11110_ (.A1(_06290_),
    .A2(\register_file[27][15] ),
    .ZN(_06294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11111_ (.A1(_06095_),
    .A2(_06293_),
    .B(_06294_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11112_ (.A1(_06290_),
    .A2(\register_file[27][16] ),
    .ZN(_06295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11113_ (.A1(_06100_),
    .A2(_06293_),
    .B(_06295_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11114_ (.A1(_06290_),
    .A2(\register_file[27][17] ),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11115_ (.A1(_06104_),
    .A2(_06293_),
    .B(_06296_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11116_ (.I(_06267_),
    .Z(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11117_ (.A1(_06297_),
    .A2(\register_file[27][18] ),
    .ZN(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11118_ (.A1(_06108_),
    .A2(_06293_),
    .B(_06298_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11119_ (.A1(_06297_),
    .A2(\register_file[27][19] ),
    .ZN(_06299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11120_ (.A1(_06113_),
    .A2(_06293_),
    .B(_06299_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11121_ (.I(_06278_),
    .Z(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11122_ (.A1(_06297_),
    .A2(\register_file[27][20] ),
    .ZN(_06301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11123_ (.A1(_06117_),
    .A2(_06300_),
    .B(_06301_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11124_ (.A1(_06297_),
    .A2(\register_file[27][21] ),
    .ZN(_06302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11125_ (.A1(_06122_),
    .A2(_06300_),
    .B(_06302_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11126_ (.A1(_06297_),
    .A2(\register_file[27][22] ),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11127_ (.A1(_06126_),
    .A2(_06300_),
    .B(_06303_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11128_ (.I(_06267_),
    .Z(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11129_ (.A1(_06304_),
    .A2(\register_file[27][23] ),
    .ZN(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11130_ (.A1(_06130_),
    .A2(_06300_),
    .B(_06305_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11131_ (.A1(_06304_),
    .A2(\register_file[27][24] ),
    .ZN(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11132_ (.A1(_06135_),
    .A2(_06300_),
    .B(_06306_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11133_ (.I(_06278_),
    .Z(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11134_ (.A1(_06304_),
    .A2(\register_file[27][25] ),
    .ZN(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11135_ (.A1(_06139_),
    .A2(_06307_),
    .B(_06308_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11136_ (.A1(_06304_),
    .A2(\register_file[27][26] ),
    .ZN(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11137_ (.A1(_06144_),
    .A2(_06307_),
    .B(_06309_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11138_ (.A1(_06304_),
    .A2(\register_file[27][27] ),
    .ZN(_06310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11139_ (.A1(_06148_),
    .A2(_06307_),
    .B(_06310_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11140_ (.A1(_06268_),
    .A2(\register_file[27][28] ),
    .ZN(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11141_ (.A1(_06152_),
    .A2(_06307_),
    .B(_06311_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11142_ (.A1(_06268_),
    .A2(\register_file[27][29] ),
    .ZN(_06312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11143_ (.A1(_06156_),
    .A2(_06307_),
    .B(_06312_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11144_ (.A1(_06268_),
    .A2(\register_file[27][30] ),
    .ZN(_06313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11145_ (.A1(_06160_),
    .A2(_06271_),
    .B(_06313_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11146_ (.A1(_06268_),
    .A2(\register_file[27][31] ),
    .ZN(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11147_ (.A1(_06164_),
    .A2(_06271_),
    .B(_06314_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11148_ (.A1(_03764_),
    .A2(net43),
    .ZN(_06315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11149_ (.I(_06315_),
    .ZN(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11150_ (.I(_06316_),
    .Z(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11151_ (.A1(_06317_),
    .A2(_04219_),
    .ZN(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11152_ (.I(_06318_),
    .Z(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11153_ (.I(_06319_),
    .Z(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11154_ (.I(_06318_),
    .Z(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11155_ (.I(_06321_),
    .Z(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11156_ (.A1(_06322_),
    .A2(\register_file[13][0] ),
    .ZN(_06323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11157_ (.A1(_06021_),
    .A2(_06320_),
    .B(_06323_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11158_ (.A1(_06322_),
    .A2(\register_file[13][1] ),
    .ZN(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11159_ (.A1(_06033_),
    .A2(_06320_),
    .B(_06324_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11160_ (.A1(_06322_),
    .A2(\register_file[13][2] ),
    .ZN(_06325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11161_ (.A1(_06037_),
    .A2(_06320_),
    .B(_06325_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11162_ (.I(_06321_),
    .Z(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11163_ (.A1(_06326_),
    .A2(\register_file[13][3] ),
    .ZN(_06327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11164_ (.A1(_06041_),
    .A2(_06320_),
    .B(_06327_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11165_ (.A1(_06326_),
    .A2(\register_file[13][4] ),
    .ZN(_06328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11166_ (.A1(_06046_),
    .A2(_06320_),
    .B(_06328_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11167_ (.I(_06321_),
    .Z(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11168_ (.I(_06329_),
    .Z(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11169_ (.A1(_06326_),
    .A2(\register_file[13][5] ),
    .ZN(_06331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11170_ (.A1(_06050_),
    .A2(_06330_),
    .B(_06331_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11171_ (.A1(_06326_),
    .A2(\register_file[13][6] ),
    .ZN(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11172_ (.A1(_06056_),
    .A2(_06330_),
    .B(_06332_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11173_ (.A1(_06326_),
    .A2(\register_file[13][7] ),
    .ZN(_06333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11174_ (.A1(_06060_),
    .A2(_06330_),
    .B(_06333_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11175_ (.I(_06321_),
    .Z(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11176_ (.A1(_06334_),
    .A2(\register_file[13][8] ),
    .ZN(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11177_ (.A1(_06064_),
    .A2(_06330_),
    .B(_06335_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11178_ (.A1(_06334_),
    .A2(\register_file[13][9] ),
    .ZN(_06336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11179_ (.A1(_06069_),
    .A2(_06330_),
    .B(_06336_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11180_ (.I(_06329_),
    .Z(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11181_ (.A1(_06334_),
    .A2(\register_file[13][10] ),
    .ZN(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11182_ (.A1(_06073_),
    .A2(_06337_),
    .B(_06338_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11183_ (.A1(_06334_),
    .A2(\register_file[13][11] ),
    .ZN(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11184_ (.A1(_06078_),
    .A2(_06337_),
    .B(_06339_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11185_ (.A1(_06334_),
    .A2(\register_file[13][12] ),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11186_ (.A1(_06082_),
    .A2(_06337_),
    .B(_06340_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11187_ (.I(_06321_),
    .Z(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11188_ (.A1(_06341_),
    .A2(\register_file[13][13] ),
    .ZN(_06342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11189_ (.A1(_06086_),
    .A2(_06337_),
    .B(_06342_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11190_ (.A1(_06341_),
    .A2(\register_file[13][14] ),
    .ZN(_06343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11191_ (.A1(_06091_),
    .A2(_06337_),
    .B(_06343_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11192_ (.I(_06329_),
    .Z(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11193_ (.A1(_06341_),
    .A2(\register_file[13][15] ),
    .ZN(_06345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11194_ (.A1(_06095_),
    .A2(_06344_),
    .B(_06345_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11195_ (.A1(_06341_),
    .A2(\register_file[13][16] ),
    .ZN(_06346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11196_ (.A1(_06100_),
    .A2(_06344_),
    .B(_06346_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11197_ (.A1(_06341_),
    .A2(\register_file[13][17] ),
    .ZN(_06347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11198_ (.A1(_06104_),
    .A2(_06344_),
    .B(_06347_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11199_ (.I(_06318_),
    .Z(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11200_ (.A1(_06348_),
    .A2(\register_file[13][18] ),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11201_ (.A1(_06108_),
    .A2(_06344_),
    .B(_06349_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11202_ (.A1(_06348_),
    .A2(\register_file[13][19] ),
    .ZN(_06350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11203_ (.A1(_06113_),
    .A2(_06344_),
    .B(_06350_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11204_ (.I(_06329_),
    .Z(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11205_ (.A1(_06348_),
    .A2(\register_file[13][20] ),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11206_ (.A1(_06117_),
    .A2(_06351_),
    .B(_06352_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11207_ (.A1(_06348_),
    .A2(\register_file[13][21] ),
    .ZN(_06353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11208_ (.A1(_06122_),
    .A2(_06351_),
    .B(_06353_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11209_ (.A1(_06348_),
    .A2(\register_file[13][22] ),
    .ZN(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11210_ (.A1(_06126_),
    .A2(_06351_),
    .B(_06354_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11211_ (.I(_06318_),
    .Z(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11212_ (.A1(_06355_),
    .A2(\register_file[13][23] ),
    .ZN(_06356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11213_ (.A1(_06130_),
    .A2(_06351_),
    .B(_06356_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11214_ (.A1(_06355_),
    .A2(\register_file[13][24] ),
    .ZN(_06357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11215_ (.A1(_06135_),
    .A2(_06351_),
    .B(_06357_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11216_ (.I(_06329_),
    .Z(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11217_ (.A1(_06355_),
    .A2(\register_file[13][25] ),
    .ZN(_06359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11218_ (.A1(_06139_),
    .A2(_06358_),
    .B(_06359_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11219_ (.A1(_06355_),
    .A2(\register_file[13][26] ),
    .ZN(_06360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11220_ (.A1(_06144_),
    .A2(_06358_),
    .B(_06360_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11221_ (.A1(_06355_),
    .A2(\register_file[13][27] ),
    .ZN(_06361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11222_ (.A1(_06148_),
    .A2(_06358_),
    .B(_06361_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11223_ (.A1(_06319_),
    .A2(\register_file[13][28] ),
    .ZN(_06362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11224_ (.A1(_06152_),
    .A2(_06358_),
    .B(_06362_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11225_ (.A1(_06319_),
    .A2(\register_file[13][29] ),
    .ZN(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11226_ (.A1(_06156_),
    .A2(_06358_),
    .B(_06363_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11227_ (.A1(_06319_),
    .A2(\register_file[13][30] ),
    .ZN(_06364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11228_ (.A1(_06160_),
    .A2(_06322_),
    .B(_06364_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11229_ (.A1(_06319_),
    .A2(\register_file[13][31] ),
    .ZN(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11230_ (.A1(_06164_),
    .A2(_06322_),
    .B(_06365_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11231_ (.I(_06020_),
    .Z(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11232_ (.A1(_06266_),
    .A2(_03855_),
    .ZN(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11233_ (.I(_06367_),
    .Z(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11234_ (.I(_06368_),
    .Z(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11235_ (.I(_06367_),
    .Z(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11236_ (.I(_06370_),
    .Z(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11237_ (.A1(_06371_),
    .A2(\register_file[19][0] ),
    .ZN(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11238_ (.A1(_06366_),
    .A2(_06369_),
    .B(_06372_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11239_ (.I(_06032_),
    .Z(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11240_ (.A1(_06371_),
    .A2(\register_file[19][1] ),
    .ZN(_06374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11241_ (.A1(_06373_),
    .A2(_06369_),
    .B(_06374_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11242_ (.I(_06036_),
    .Z(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11243_ (.A1(_06371_),
    .A2(\register_file[19][2] ),
    .ZN(_06376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11244_ (.A1(_06375_),
    .A2(_06369_),
    .B(_06376_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11245_ (.I(_06040_),
    .Z(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11246_ (.I(_06370_),
    .Z(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11247_ (.A1(_06378_),
    .A2(\register_file[19][3] ),
    .ZN(_06379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11248_ (.A1(_06377_),
    .A2(_06369_),
    .B(_06379_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11249_ (.I(_06045_),
    .Z(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11250_ (.A1(_06378_),
    .A2(\register_file[19][4] ),
    .ZN(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11251_ (.A1(_06380_),
    .A2(_06369_),
    .B(_06381_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11252_ (.I(_06049_),
    .Z(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11253_ (.I(_06370_),
    .Z(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11254_ (.I(_06383_),
    .Z(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11255_ (.A1(_06378_),
    .A2(\register_file[19][5] ),
    .ZN(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11256_ (.A1(_06382_),
    .A2(_06384_),
    .B(_06385_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11257_ (.I(_06055_),
    .Z(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11258_ (.A1(_06378_),
    .A2(\register_file[19][6] ),
    .ZN(_06387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11259_ (.A1(_06386_),
    .A2(_06384_),
    .B(_06387_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11260_ (.I(_06059_),
    .Z(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11261_ (.A1(_06378_),
    .A2(\register_file[19][7] ),
    .ZN(_06389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11262_ (.A1(_06388_),
    .A2(_06384_),
    .B(_06389_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11263_ (.I(_06063_),
    .Z(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11264_ (.I(_06370_),
    .Z(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11265_ (.A1(_06391_),
    .A2(\register_file[19][8] ),
    .ZN(_06392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11266_ (.A1(_06390_),
    .A2(_06384_),
    .B(_06392_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11267_ (.I(_06068_),
    .Z(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11268_ (.A1(_06391_),
    .A2(\register_file[19][9] ),
    .ZN(_06394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11269_ (.A1(_06393_),
    .A2(_06384_),
    .B(_06394_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11270_ (.I(_06072_),
    .Z(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11271_ (.I(_06383_),
    .Z(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11272_ (.A1(_06391_),
    .A2(\register_file[19][10] ),
    .ZN(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11273_ (.A1(_06395_),
    .A2(_06396_),
    .B(_06397_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11274_ (.I(_06077_),
    .Z(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11275_ (.A1(_06391_),
    .A2(\register_file[19][11] ),
    .ZN(_06399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11276_ (.A1(_06398_),
    .A2(_06396_),
    .B(_06399_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11277_ (.I(_06081_),
    .Z(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11278_ (.A1(_06391_),
    .A2(\register_file[19][12] ),
    .ZN(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11279_ (.A1(_06400_),
    .A2(_06396_),
    .B(_06401_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11280_ (.I(_06085_),
    .Z(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11281_ (.I(_06370_),
    .Z(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11282_ (.A1(_06403_),
    .A2(\register_file[19][13] ),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11283_ (.A1(_06402_),
    .A2(_06396_),
    .B(_06404_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11284_ (.I(_06090_),
    .Z(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11285_ (.A1(_06403_),
    .A2(\register_file[19][14] ),
    .ZN(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11286_ (.A1(_06405_),
    .A2(_06396_),
    .B(_06406_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11287_ (.I(_06094_),
    .Z(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11288_ (.I(_06383_),
    .Z(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11289_ (.A1(_06403_),
    .A2(\register_file[19][15] ),
    .ZN(_06409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11290_ (.A1(_06407_),
    .A2(_06408_),
    .B(_06409_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11291_ (.I(_06099_),
    .Z(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11292_ (.A1(_06403_),
    .A2(\register_file[19][16] ),
    .ZN(_06411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11293_ (.A1(_06410_),
    .A2(_06408_),
    .B(_06411_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11294_ (.I(_06103_),
    .Z(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11295_ (.A1(_06403_),
    .A2(\register_file[19][17] ),
    .ZN(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11296_ (.A1(_06412_),
    .A2(_06408_),
    .B(_06413_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11297_ (.I(_06107_),
    .Z(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11298_ (.I(_06367_),
    .Z(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11299_ (.A1(_06415_),
    .A2(\register_file[19][18] ),
    .ZN(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11300_ (.A1(_06414_),
    .A2(_06408_),
    .B(_06416_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11301_ (.I(_06112_),
    .Z(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11302_ (.A1(_06415_),
    .A2(\register_file[19][19] ),
    .ZN(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11303_ (.A1(_06417_),
    .A2(_06408_),
    .B(_06418_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11304_ (.I(_06116_),
    .Z(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11305_ (.I(_06383_),
    .Z(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11306_ (.A1(_06415_),
    .A2(\register_file[19][20] ),
    .ZN(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11307_ (.A1(_06419_),
    .A2(_06420_),
    .B(_06421_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11308_ (.I(_06121_),
    .Z(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11309_ (.A1(_06415_),
    .A2(\register_file[19][21] ),
    .ZN(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11310_ (.A1(_06422_),
    .A2(_06420_),
    .B(_06423_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11311_ (.I(_06125_),
    .Z(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11312_ (.A1(_06415_),
    .A2(\register_file[19][22] ),
    .ZN(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11313_ (.A1(_06424_),
    .A2(_06420_),
    .B(_06425_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11314_ (.I(_06129_),
    .Z(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11315_ (.I(_06367_),
    .Z(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11316_ (.A1(_06427_),
    .A2(\register_file[19][23] ),
    .ZN(_06428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11317_ (.A1(_06426_),
    .A2(_06420_),
    .B(_06428_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11318_ (.I(_06134_),
    .Z(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11319_ (.A1(_06427_),
    .A2(\register_file[19][24] ),
    .ZN(_06430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11320_ (.A1(_06429_),
    .A2(_06420_),
    .B(_06430_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11321_ (.I(_06138_),
    .Z(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11322_ (.I(_06383_),
    .Z(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11323_ (.A1(_06427_),
    .A2(\register_file[19][25] ),
    .ZN(_06433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11324_ (.A1(_06431_),
    .A2(_06432_),
    .B(_06433_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11325_ (.I(_06143_),
    .Z(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11326_ (.A1(_06427_),
    .A2(\register_file[19][26] ),
    .ZN(_06435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11327_ (.A1(_06434_),
    .A2(_06432_),
    .B(_06435_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11328_ (.I(_06147_),
    .Z(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11329_ (.A1(_06427_),
    .A2(\register_file[19][27] ),
    .ZN(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11330_ (.A1(_06436_),
    .A2(_06432_),
    .B(_06437_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11331_ (.I(_06151_),
    .Z(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11332_ (.A1(_06368_),
    .A2(\register_file[19][28] ),
    .ZN(_06439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11333_ (.A1(_06438_),
    .A2(_06432_),
    .B(_06439_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11334_ (.I(_06155_),
    .Z(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11335_ (.A1(_06368_),
    .A2(\register_file[19][29] ),
    .ZN(_06441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11336_ (.A1(_06440_),
    .A2(_06432_),
    .B(_06441_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11337_ (.I(_06159_),
    .Z(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11338_ (.A1(_06368_),
    .A2(\register_file[19][30] ),
    .ZN(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11339_ (.A1(_06442_),
    .A2(_06371_),
    .B(_06443_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11340_ (.I(_06163_),
    .Z(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11341_ (.A1(_06368_),
    .A2(\register_file[19][31] ),
    .ZN(_06445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11342_ (.A1(_06444_),
    .A2(_06371_),
    .B(_06445_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11343_ (.A1(_06024_),
    .A2(_03794_),
    .ZN(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11344_ (.I(_06446_),
    .Z(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11345_ (.I(_06447_),
    .Z(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11346_ (.I(_06446_),
    .Z(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11347_ (.I(_06449_),
    .Z(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11348_ (.A1(_06450_),
    .A2(\register_file[26][0] ),
    .ZN(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11349_ (.A1(_06366_),
    .A2(_06448_),
    .B(_06451_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11350_ (.A1(_06450_),
    .A2(\register_file[26][1] ),
    .ZN(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11351_ (.A1(_06373_),
    .A2(_06448_),
    .B(_06452_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11352_ (.A1(_06450_),
    .A2(\register_file[26][2] ),
    .ZN(_06453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11353_ (.A1(_06375_),
    .A2(_06448_),
    .B(_06453_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11354_ (.I(_06449_),
    .Z(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11355_ (.A1(_06454_),
    .A2(\register_file[26][3] ),
    .ZN(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11356_ (.A1(_06377_),
    .A2(_06448_),
    .B(_06455_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11357_ (.A1(_06454_),
    .A2(\register_file[26][4] ),
    .ZN(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11358_ (.A1(_06380_),
    .A2(_06448_),
    .B(_06456_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11359_ (.I(_06449_),
    .Z(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11360_ (.I(_06457_),
    .Z(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11361_ (.A1(_06454_),
    .A2(\register_file[26][5] ),
    .ZN(_06459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11362_ (.A1(_06382_),
    .A2(_06458_),
    .B(_06459_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11363_ (.A1(_06454_),
    .A2(\register_file[26][6] ),
    .ZN(_06460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11364_ (.A1(_06386_),
    .A2(_06458_),
    .B(_06460_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11365_ (.A1(_06454_),
    .A2(\register_file[26][7] ),
    .ZN(_06461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11366_ (.A1(_06388_),
    .A2(_06458_),
    .B(_06461_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11367_ (.I(_06449_),
    .Z(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11368_ (.A1(_06462_),
    .A2(\register_file[26][8] ),
    .ZN(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11369_ (.A1(_06390_),
    .A2(_06458_),
    .B(_06463_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11370_ (.A1(_06462_),
    .A2(\register_file[26][9] ),
    .ZN(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11371_ (.A1(_06393_),
    .A2(_06458_),
    .B(_06464_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11372_ (.I(_06457_),
    .Z(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11373_ (.A1(_06462_),
    .A2(\register_file[26][10] ),
    .ZN(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11374_ (.A1(_06395_),
    .A2(_06465_),
    .B(_06466_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11375_ (.A1(_06462_),
    .A2(\register_file[26][11] ),
    .ZN(_06467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11376_ (.A1(_06398_),
    .A2(_06465_),
    .B(_06467_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11377_ (.A1(_06462_),
    .A2(\register_file[26][12] ),
    .ZN(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11378_ (.A1(_06400_),
    .A2(_06465_),
    .B(_06468_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11379_ (.I(_06449_),
    .Z(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11380_ (.A1(_06469_),
    .A2(\register_file[26][13] ),
    .ZN(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11381_ (.A1(_06402_),
    .A2(_06465_),
    .B(_06470_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11382_ (.A1(_06469_),
    .A2(\register_file[26][14] ),
    .ZN(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11383_ (.A1(_06405_),
    .A2(_06465_),
    .B(_06471_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11384_ (.I(_06457_),
    .Z(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11385_ (.A1(_06469_),
    .A2(\register_file[26][15] ),
    .ZN(_06473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11386_ (.A1(_06407_),
    .A2(_06472_),
    .B(_06473_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11387_ (.A1(_06469_),
    .A2(\register_file[26][16] ),
    .ZN(_06474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11388_ (.A1(_06410_),
    .A2(_06472_),
    .B(_06474_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11389_ (.A1(_06469_),
    .A2(\register_file[26][17] ),
    .ZN(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11390_ (.A1(_06412_),
    .A2(_06472_),
    .B(_06475_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11391_ (.I(_06446_),
    .Z(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11392_ (.A1(_06476_),
    .A2(\register_file[26][18] ),
    .ZN(_06477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11393_ (.A1(_06414_),
    .A2(_06472_),
    .B(_06477_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11394_ (.A1(_06476_),
    .A2(\register_file[26][19] ),
    .ZN(_06478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11395_ (.A1(_06417_),
    .A2(_06472_),
    .B(_06478_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11396_ (.I(_06457_),
    .Z(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11397_ (.A1(_06476_),
    .A2(\register_file[26][20] ),
    .ZN(_06480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11398_ (.A1(_06419_),
    .A2(_06479_),
    .B(_06480_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11399_ (.A1(_06476_),
    .A2(\register_file[26][21] ),
    .ZN(_06481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11400_ (.A1(_06422_),
    .A2(_06479_),
    .B(_06481_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11401_ (.A1(_06476_),
    .A2(\register_file[26][22] ),
    .ZN(_06482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11402_ (.A1(_06424_),
    .A2(_06479_),
    .B(_06482_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11403_ (.I(_06446_),
    .Z(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11404_ (.A1(_06483_),
    .A2(\register_file[26][23] ),
    .ZN(_06484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11405_ (.A1(_06426_),
    .A2(_06479_),
    .B(_06484_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11406_ (.A1(_06483_),
    .A2(\register_file[26][24] ),
    .ZN(_06485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11407_ (.A1(_06429_),
    .A2(_06479_),
    .B(_06485_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11408_ (.I(_06457_),
    .Z(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11409_ (.A1(_06483_),
    .A2(\register_file[26][25] ),
    .ZN(_06487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11410_ (.A1(_06431_),
    .A2(_06486_),
    .B(_06487_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11411_ (.A1(_06483_),
    .A2(\register_file[26][26] ),
    .ZN(_06488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11412_ (.A1(_06434_),
    .A2(_06486_),
    .B(_06488_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11413_ (.A1(_06483_),
    .A2(\register_file[26][27] ),
    .ZN(_06489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11414_ (.A1(_06436_),
    .A2(_06486_),
    .B(_06489_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11415_ (.A1(_06447_),
    .A2(\register_file[26][28] ),
    .ZN(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11416_ (.A1(_06438_),
    .A2(_06486_),
    .B(_06490_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11417_ (.A1(_06447_),
    .A2(\register_file[26][29] ),
    .ZN(_06491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11418_ (.A1(_06440_),
    .A2(_06486_),
    .B(_06491_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11419_ (.A1(_06447_),
    .A2(\register_file[26][30] ),
    .ZN(_06492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11420_ (.A1(_06442_),
    .A2(_06450_),
    .B(_06492_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11421_ (.A1(_06447_),
    .A2(\register_file[26][31] ),
    .ZN(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11422_ (.A1(_06444_),
    .A2(_06450_),
    .B(_06493_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11423_ (.A1(_06216_),
    .A2(_04219_),
    .ZN(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11424_ (.I(_06494_),
    .Z(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11425_ (.I(_06495_),
    .Z(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11426_ (.I(_06494_),
    .Z(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11427_ (.I(_06497_),
    .Z(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11428_ (.A1(_06498_),
    .A2(\register_file[12][0] ),
    .ZN(_06499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11429_ (.A1(_06366_),
    .A2(_06496_),
    .B(_06499_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11430_ (.A1(_06498_),
    .A2(\register_file[12][1] ),
    .ZN(_06500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11431_ (.A1(_06373_),
    .A2(_06496_),
    .B(_06500_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11432_ (.A1(_06498_),
    .A2(\register_file[12][2] ),
    .ZN(_06501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11433_ (.A1(_06375_),
    .A2(_06496_),
    .B(_06501_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11434_ (.I(_06497_),
    .Z(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11435_ (.A1(_06502_),
    .A2(\register_file[12][3] ),
    .ZN(_06503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11436_ (.A1(_06377_),
    .A2(_06496_),
    .B(_06503_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11437_ (.A1(_06502_),
    .A2(\register_file[12][4] ),
    .ZN(_06504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11438_ (.A1(_06380_),
    .A2(_06496_),
    .B(_06504_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11439_ (.I(_06497_),
    .Z(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11440_ (.I(_06505_),
    .Z(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11441_ (.A1(_06502_),
    .A2(\register_file[12][5] ),
    .ZN(_06507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11442_ (.A1(_06382_),
    .A2(_06506_),
    .B(_06507_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11443_ (.A1(_06502_),
    .A2(\register_file[12][6] ),
    .ZN(_06508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11444_ (.A1(_06386_),
    .A2(_06506_),
    .B(_06508_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11445_ (.A1(_06502_),
    .A2(\register_file[12][7] ),
    .ZN(_06509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11446_ (.A1(_06388_),
    .A2(_06506_),
    .B(_06509_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11447_ (.I(_06497_),
    .Z(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11448_ (.A1(_06510_),
    .A2(\register_file[12][8] ),
    .ZN(_06511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11449_ (.A1(_06390_),
    .A2(_06506_),
    .B(_06511_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11450_ (.A1(_06510_),
    .A2(\register_file[12][9] ),
    .ZN(_06512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11451_ (.A1(_06393_),
    .A2(_06506_),
    .B(_06512_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11452_ (.I(_06505_),
    .Z(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11453_ (.A1(_06510_),
    .A2(\register_file[12][10] ),
    .ZN(_06514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11454_ (.A1(_06395_),
    .A2(_06513_),
    .B(_06514_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11455_ (.A1(_06510_),
    .A2(\register_file[12][11] ),
    .ZN(_06515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11456_ (.A1(_06398_),
    .A2(_06513_),
    .B(_06515_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11457_ (.A1(_06510_),
    .A2(\register_file[12][12] ),
    .ZN(_06516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11458_ (.A1(_06400_),
    .A2(_06513_),
    .B(_06516_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11459_ (.I(_06497_),
    .Z(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11460_ (.A1(_06517_),
    .A2(\register_file[12][13] ),
    .ZN(_06518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11461_ (.A1(_06402_),
    .A2(_06513_),
    .B(_06518_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11462_ (.A1(_06517_),
    .A2(\register_file[12][14] ),
    .ZN(_06519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11463_ (.A1(_06405_),
    .A2(_06513_),
    .B(_06519_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11464_ (.I(_06505_),
    .Z(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11465_ (.A1(_06517_),
    .A2(\register_file[12][15] ),
    .ZN(_06521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11466_ (.A1(_06407_),
    .A2(_06520_),
    .B(_06521_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11467_ (.A1(_06517_),
    .A2(\register_file[12][16] ),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11468_ (.A1(_06410_),
    .A2(_06520_),
    .B(_06522_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11469_ (.A1(_06517_),
    .A2(\register_file[12][17] ),
    .ZN(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11470_ (.A1(_06412_),
    .A2(_06520_),
    .B(_06523_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11471_ (.I(_06494_),
    .Z(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11472_ (.A1(_06524_),
    .A2(\register_file[12][18] ),
    .ZN(_06525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11473_ (.A1(_06414_),
    .A2(_06520_),
    .B(_06525_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11474_ (.A1(_06524_),
    .A2(\register_file[12][19] ),
    .ZN(_06526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11475_ (.A1(_06417_),
    .A2(_06520_),
    .B(_06526_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11476_ (.I(_06505_),
    .Z(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11477_ (.A1(_06524_),
    .A2(\register_file[12][20] ),
    .ZN(_06528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11478_ (.A1(_06419_),
    .A2(_06527_),
    .B(_06528_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11479_ (.A1(_06524_),
    .A2(\register_file[12][21] ),
    .ZN(_06529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11480_ (.A1(_06422_),
    .A2(_06527_),
    .B(_06529_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11481_ (.A1(_06524_),
    .A2(\register_file[12][22] ),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11482_ (.A1(_06424_),
    .A2(_06527_),
    .B(_06530_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11483_ (.I(_06494_),
    .Z(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11484_ (.A1(_06531_),
    .A2(\register_file[12][23] ),
    .ZN(_06532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11485_ (.A1(_06426_),
    .A2(_06527_),
    .B(_06532_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11486_ (.A1(_06531_),
    .A2(\register_file[12][24] ),
    .ZN(_06533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11487_ (.A1(_06429_),
    .A2(_06527_),
    .B(_06533_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11488_ (.I(_06505_),
    .Z(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11489_ (.A1(_06531_),
    .A2(\register_file[12][25] ),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11490_ (.A1(_06431_),
    .A2(_06534_),
    .B(_06535_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11491_ (.A1(_06531_),
    .A2(\register_file[12][26] ),
    .ZN(_06536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11492_ (.A1(_06434_),
    .A2(_06534_),
    .B(_06536_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11493_ (.A1(_06531_),
    .A2(\register_file[12][27] ),
    .ZN(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11494_ (.A1(_06436_),
    .A2(_06534_),
    .B(_06537_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11495_ (.A1(_06495_),
    .A2(\register_file[12][28] ),
    .ZN(_06538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11496_ (.A1(_06438_),
    .A2(_06534_),
    .B(_06538_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11497_ (.A1(_06495_),
    .A2(\register_file[12][29] ),
    .ZN(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11498_ (.A1(_06440_),
    .A2(_06534_),
    .B(_06539_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11499_ (.A1(_06495_),
    .A2(\register_file[12][30] ),
    .ZN(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11500_ (.A1(_06442_),
    .A2(_06498_),
    .B(_06540_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11501_ (.A1(_06495_),
    .A2(\register_file[12][31] ),
    .ZN(_06541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11502_ (.A1(_06444_),
    .A2(_06498_),
    .B(_06541_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11503_ (.A1(_06266_),
    .A2(_04001_),
    .ZN(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11504_ (.I(_06542_),
    .Z(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11505_ (.I(_06543_),
    .Z(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11506_ (.I(_06542_),
    .Z(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11507_ (.I(_06545_),
    .Z(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11508_ (.A1(_06546_),
    .A2(\register_file[11][0] ),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11509_ (.A1(_06366_),
    .A2(_06544_),
    .B(_06547_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11510_ (.A1(_06546_),
    .A2(\register_file[11][1] ),
    .ZN(_06548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11511_ (.A1(_06373_),
    .A2(_06544_),
    .B(_06548_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11512_ (.A1(_06546_),
    .A2(\register_file[11][2] ),
    .ZN(_06549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11513_ (.A1(_06375_),
    .A2(_06544_),
    .B(_06549_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11514_ (.I(_06545_),
    .Z(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11515_ (.A1(_06550_),
    .A2(\register_file[11][3] ),
    .ZN(_06551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11516_ (.A1(_06377_),
    .A2(_06544_),
    .B(_06551_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11517_ (.A1(_06550_),
    .A2(\register_file[11][4] ),
    .ZN(_06552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11518_ (.A1(_06380_),
    .A2(_06544_),
    .B(_06552_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11519_ (.I(_06545_),
    .Z(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11520_ (.I(_06553_),
    .Z(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11521_ (.A1(_06550_),
    .A2(\register_file[11][5] ),
    .ZN(_06555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11522_ (.A1(_06382_),
    .A2(_06554_),
    .B(_06555_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11523_ (.A1(_06550_),
    .A2(\register_file[11][6] ),
    .ZN(_06556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11524_ (.A1(_06386_),
    .A2(_06554_),
    .B(_06556_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11525_ (.A1(_06550_),
    .A2(\register_file[11][7] ),
    .ZN(_06557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11526_ (.A1(_06388_),
    .A2(_06554_),
    .B(_06557_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11527_ (.I(_06545_),
    .Z(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11528_ (.A1(_06558_),
    .A2(\register_file[11][8] ),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11529_ (.A1(_06390_),
    .A2(_06554_),
    .B(_06559_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11530_ (.A1(_06558_),
    .A2(\register_file[11][9] ),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11531_ (.A1(_06393_),
    .A2(_06554_),
    .B(_06560_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11532_ (.I(_06553_),
    .Z(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11533_ (.A1(_06558_),
    .A2(\register_file[11][10] ),
    .ZN(_06562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11534_ (.A1(_06395_),
    .A2(_06561_),
    .B(_06562_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11535_ (.A1(_06558_),
    .A2(\register_file[11][11] ),
    .ZN(_06563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11536_ (.A1(_06398_),
    .A2(_06561_),
    .B(_06563_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11537_ (.A1(_06558_),
    .A2(\register_file[11][12] ),
    .ZN(_06564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11538_ (.A1(_06400_),
    .A2(_06561_),
    .B(_06564_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11539_ (.I(_06545_),
    .Z(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11540_ (.A1(_06565_),
    .A2(\register_file[11][13] ),
    .ZN(_06566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11541_ (.A1(_06402_),
    .A2(_06561_),
    .B(_06566_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11542_ (.A1(_06565_),
    .A2(\register_file[11][14] ),
    .ZN(_06567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11543_ (.A1(_06405_),
    .A2(_06561_),
    .B(_06567_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11544_ (.I(_06553_),
    .Z(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11545_ (.A1(_06565_),
    .A2(\register_file[11][15] ),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11546_ (.A1(_06407_),
    .A2(_06568_),
    .B(_06569_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11547_ (.A1(_06565_),
    .A2(\register_file[11][16] ),
    .ZN(_06570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11548_ (.A1(_06410_),
    .A2(_06568_),
    .B(_06570_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11549_ (.A1(_06565_),
    .A2(\register_file[11][17] ),
    .ZN(_06571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11550_ (.A1(_06412_),
    .A2(_06568_),
    .B(_06571_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11551_ (.I(_06542_),
    .Z(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11552_ (.A1(_06572_),
    .A2(\register_file[11][18] ),
    .ZN(_06573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11553_ (.A1(_06414_),
    .A2(_06568_),
    .B(_06573_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11554_ (.A1(_06572_),
    .A2(\register_file[11][19] ),
    .ZN(_06574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11555_ (.A1(_06417_),
    .A2(_06568_),
    .B(_06574_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11556_ (.I(_06553_),
    .Z(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11557_ (.A1(_06572_),
    .A2(\register_file[11][20] ),
    .ZN(_06576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11558_ (.A1(_06419_),
    .A2(_06575_),
    .B(_06576_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11559_ (.A1(_06572_),
    .A2(\register_file[11][21] ),
    .ZN(_06577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11560_ (.A1(_06422_),
    .A2(_06575_),
    .B(_06577_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11561_ (.A1(_06572_),
    .A2(\register_file[11][22] ),
    .ZN(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11562_ (.A1(_06424_),
    .A2(_06575_),
    .B(_06578_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11563_ (.I(_06542_),
    .Z(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11564_ (.A1(_06579_),
    .A2(\register_file[11][23] ),
    .ZN(_06580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11565_ (.A1(_06426_),
    .A2(_06575_),
    .B(_06580_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11566_ (.A1(_06579_),
    .A2(\register_file[11][24] ),
    .ZN(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11567_ (.A1(_06429_),
    .A2(_06575_),
    .B(_06581_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11568_ (.I(_06553_),
    .Z(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11569_ (.A1(_06579_),
    .A2(\register_file[11][25] ),
    .ZN(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11570_ (.A1(_06431_),
    .A2(_06582_),
    .B(_06583_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11571_ (.A1(_06579_),
    .A2(\register_file[11][26] ),
    .ZN(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11572_ (.A1(_06434_),
    .A2(_06582_),
    .B(_06584_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11573_ (.A1(_06579_),
    .A2(\register_file[11][27] ),
    .ZN(_06585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11574_ (.A1(_06436_),
    .A2(_06582_),
    .B(_06585_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11575_ (.A1(_06543_),
    .A2(\register_file[11][28] ),
    .ZN(_06586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11576_ (.A1(_06438_),
    .A2(_06582_),
    .B(_06586_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11577_ (.A1(_06543_),
    .A2(\register_file[11][29] ),
    .ZN(_06587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11578_ (.A1(_06440_),
    .A2(_06582_),
    .B(_06587_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11579_ (.A1(_06543_),
    .A2(\register_file[11][30] ),
    .ZN(_06588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11580_ (.A1(_06442_),
    .A2(_06546_),
    .B(_06588_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11581_ (.A1(_06543_),
    .A2(\register_file[11][31] ),
    .ZN(_06589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11582_ (.A1(_06444_),
    .A2(_06546_),
    .B(_06589_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11583_ (.A1(_06024_),
    .A2(_04001_),
    .ZN(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11584_ (.I(_06590_),
    .Z(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11585_ (.I(_06591_),
    .Z(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11586_ (.I(_06590_),
    .Z(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11587_ (.I(_06593_),
    .Z(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11588_ (.A1(_06594_),
    .A2(\register_file[10][0] ),
    .ZN(_06595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11589_ (.A1(_06366_),
    .A2(_06592_),
    .B(_06595_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11590_ (.A1(_06594_),
    .A2(\register_file[10][1] ),
    .ZN(_06596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11591_ (.A1(_06373_),
    .A2(_06592_),
    .B(_06596_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11592_ (.A1(_06594_),
    .A2(\register_file[10][2] ),
    .ZN(_06597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11593_ (.A1(_06375_),
    .A2(_06592_),
    .B(_06597_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11594_ (.I(_06593_),
    .Z(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11595_ (.A1(_06598_),
    .A2(\register_file[10][3] ),
    .ZN(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11596_ (.A1(_06377_),
    .A2(_06592_),
    .B(_06599_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11597_ (.A1(_06598_),
    .A2(\register_file[10][4] ),
    .ZN(_06600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11598_ (.A1(_06380_),
    .A2(_06592_),
    .B(_06600_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11599_ (.I(_06593_),
    .Z(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11600_ (.I(_06601_),
    .Z(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11601_ (.A1(_06598_),
    .A2(\register_file[10][5] ),
    .ZN(_06603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11602_ (.A1(_06382_),
    .A2(_06602_),
    .B(_06603_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11603_ (.A1(_06598_),
    .A2(\register_file[10][6] ),
    .ZN(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11604_ (.A1(_06386_),
    .A2(_06602_),
    .B(_06604_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11605_ (.A1(_06598_),
    .A2(\register_file[10][7] ),
    .ZN(_06605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11606_ (.A1(_06388_),
    .A2(_06602_),
    .B(_06605_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11607_ (.I(_06593_),
    .Z(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11608_ (.A1(_06606_),
    .A2(\register_file[10][8] ),
    .ZN(_06607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11609_ (.A1(_06390_),
    .A2(_06602_),
    .B(_06607_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11610_ (.A1(_06606_),
    .A2(\register_file[10][9] ),
    .ZN(_06608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11611_ (.A1(_06393_),
    .A2(_06602_),
    .B(_06608_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11612_ (.I(_06601_),
    .Z(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11613_ (.A1(_06606_),
    .A2(\register_file[10][10] ),
    .ZN(_06610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11614_ (.A1(_06395_),
    .A2(_06609_),
    .B(_06610_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11615_ (.A1(_06606_),
    .A2(\register_file[10][11] ),
    .ZN(_06611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11616_ (.A1(_06398_),
    .A2(_06609_),
    .B(_06611_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11617_ (.A1(_06606_),
    .A2(\register_file[10][12] ),
    .ZN(_06612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11618_ (.A1(_06400_),
    .A2(_06609_),
    .B(_06612_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11619_ (.I(_06593_),
    .Z(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11620_ (.A1(_06613_),
    .A2(\register_file[10][13] ),
    .ZN(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11621_ (.A1(_06402_),
    .A2(_06609_),
    .B(_06614_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11622_ (.A1(_06613_),
    .A2(\register_file[10][14] ),
    .ZN(_06615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11623_ (.A1(_06405_),
    .A2(_06609_),
    .B(_06615_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11624_ (.I(_06601_),
    .Z(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11625_ (.A1(_06613_),
    .A2(\register_file[10][15] ),
    .ZN(_06617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11626_ (.A1(_06407_),
    .A2(_06616_),
    .B(_06617_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11627_ (.A1(_06613_),
    .A2(\register_file[10][16] ),
    .ZN(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11628_ (.A1(_06410_),
    .A2(_06616_),
    .B(_06618_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11629_ (.A1(_06613_),
    .A2(\register_file[10][17] ),
    .ZN(_06619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11630_ (.A1(_06412_),
    .A2(_06616_),
    .B(_06619_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11631_ (.I(_06590_),
    .Z(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11632_ (.A1(_06620_),
    .A2(\register_file[10][18] ),
    .ZN(_06621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11633_ (.A1(_06414_),
    .A2(_06616_),
    .B(_06621_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11634_ (.A1(_06620_),
    .A2(\register_file[10][19] ),
    .ZN(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11635_ (.A1(_06417_),
    .A2(_06616_),
    .B(_06622_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11636_ (.I(_06601_),
    .Z(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11637_ (.A1(_06620_),
    .A2(\register_file[10][20] ),
    .ZN(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11638_ (.A1(_06419_),
    .A2(_06623_),
    .B(_06624_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11639_ (.A1(_06620_),
    .A2(\register_file[10][21] ),
    .ZN(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11640_ (.A1(_06422_),
    .A2(_06623_),
    .B(_06625_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11641_ (.A1(_06620_),
    .A2(\register_file[10][22] ),
    .ZN(_06626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11642_ (.A1(_06424_),
    .A2(_06623_),
    .B(_06626_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11643_ (.I(_06590_),
    .Z(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11644_ (.A1(_06627_),
    .A2(\register_file[10][23] ),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11645_ (.A1(_06426_),
    .A2(_06623_),
    .B(_06628_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11646_ (.A1(_06627_),
    .A2(\register_file[10][24] ),
    .ZN(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11647_ (.A1(_06429_),
    .A2(_06623_),
    .B(_06629_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11648_ (.I(_06601_),
    .Z(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11649_ (.A1(_06627_),
    .A2(\register_file[10][25] ),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11650_ (.A1(_06431_),
    .A2(_06630_),
    .B(_06631_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11651_ (.A1(_06627_),
    .A2(\register_file[10][26] ),
    .ZN(_06632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11652_ (.A1(_06434_),
    .A2(_06630_),
    .B(_06632_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11653_ (.A1(_06627_),
    .A2(\register_file[10][27] ),
    .ZN(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11654_ (.A1(_06436_),
    .A2(_06630_),
    .B(_06633_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11655_ (.A1(_06591_),
    .A2(\register_file[10][28] ),
    .ZN(_06634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11656_ (.A1(_06438_),
    .A2(_06630_),
    .B(_06634_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11657_ (.A1(_06591_),
    .A2(\register_file[10][29] ),
    .ZN(_06635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11658_ (.A1(_06440_),
    .A2(_06630_),
    .B(_06635_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11659_ (.A1(_06591_),
    .A2(\register_file[10][30] ),
    .ZN(_06636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11660_ (.A1(_06442_),
    .A2(_06594_),
    .B(_06636_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11661_ (.A1(_06591_),
    .A2(\register_file[10][31] ),
    .ZN(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11662_ (.A1(_06444_),
    .A2(_06594_),
    .B(_06637_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11663_ (.I(_06020_),
    .Z(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11664_ (.A1(_06216_),
    .A2(_03893_),
    .ZN(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11665_ (.I(_06639_),
    .Z(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11666_ (.I(_06640_),
    .Z(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11667_ (.I(_06639_),
    .Z(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11668_ (.I(_06642_),
    .Z(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11669_ (.A1(_06643_),
    .A2(\register_file[8][0] ),
    .ZN(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11670_ (.A1(_06638_),
    .A2(_06641_),
    .B(_06644_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11671_ (.I(_06032_),
    .Z(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11672_ (.A1(_06643_),
    .A2(\register_file[8][1] ),
    .ZN(_06646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11673_ (.A1(_06645_),
    .A2(_06641_),
    .B(_06646_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11674_ (.I(_06036_),
    .Z(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11675_ (.A1(_06643_),
    .A2(\register_file[8][2] ),
    .ZN(_06648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11676_ (.A1(_06647_),
    .A2(_06641_),
    .B(_06648_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11677_ (.I(_06040_),
    .Z(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11678_ (.I(_06642_),
    .Z(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11679_ (.A1(_06650_),
    .A2(\register_file[8][3] ),
    .ZN(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11680_ (.A1(_06649_),
    .A2(_06641_),
    .B(_06651_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11681_ (.I(_06045_),
    .Z(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11682_ (.A1(_06650_),
    .A2(\register_file[8][4] ),
    .ZN(_06653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11683_ (.A1(_06652_),
    .A2(_06641_),
    .B(_06653_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11684_ (.I(_06049_),
    .Z(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11685_ (.I(_06642_),
    .Z(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11686_ (.I(_06655_),
    .Z(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11687_ (.A1(_06650_),
    .A2(\register_file[8][5] ),
    .ZN(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11688_ (.A1(_06654_),
    .A2(_06656_),
    .B(_06657_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11689_ (.I(_06055_),
    .Z(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11690_ (.A1(_06650_),
    .A2(\register_file[8][6] ),
    .ZN(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11691_ (.A1(_06658_),
    .A2(_06656_),
    .B(_06659_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11692_ (.I(_06059_),
    .Z(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11693_ (.A1(_06650_),
    .A2(\register_file[8][7] ),
    .ZN(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11694_ (.A1(_06660_),
    .A2(_06656_),
    .B(_06661_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11695_ (.I(_06063_),
    .Z(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11696_ (.I(_06642_),
    .Z(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11697_ (.A1(_06663_),
    .A2(\register_file[8][8] ),
    .ZN(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11698_ (.A1(_06662_),
    .A2(_06656_),
    .B(_06664_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11699_ (.I(_06068_),
    .Z(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11700_ (.A1(_06663_),
    .A2(\register_file[8][9] ),
    .ZN(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11701_ (.A1(_06665_),
    .A2(_06656_),
    .B(_06666_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11702_ (.I(_06072_),
    .Z(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11703_ (.I(_06655_),
    .Z(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11704_ (.A1(_06663_),
    .A2(\register_file[8][10] ),
    .ZN(_06669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11705_ (.A1(_06667_),
    .A2(_06668_),
    .B(_06669_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11706_ (.I(_06077_),
    .Z(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11707_ (.A1(_06663_),
    .A2(\register_file[8][11] ),
    .ZN(_06671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11708_ (.A1(_06670_),
    .A2(_06668_),
    .B(_06671_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11709_ (.I(_06081_),
    .Z(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11710_ (.A1(_06663_),
    .A2(\register_file[8][12] ),
    .ZN(_06673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11711_ (.A1(_06672_),
    .A2(_06668_),
    .B(_06673_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11712_ (.I(_06085_),
    .Z(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11713_ (.I(_06642_),
    .Z(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11714_ (.A1(_06675_),
    .A2(\register_file[8][13] ),
    .ZN(_06676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11715_ (.A1(_06674_),
    .A2(_06668_),
    .B(_06676_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11716_ (.I(_06090_),
    .Z(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11717_ (.A1(_06675_),
    .A2(\register_file[8][14] ),
    .ZN(_06678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11718_ (.A1(_06677_),
    .A2(_06668_),
    .B(_06678_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11719_ (.I(_06094_),
    .Z(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11720_ (.I(_06655_),
    .Z(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11721_ (.A1(_06675_),
    .A2(\register_file[8][15] ),
    .ZN(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11722_ (.A1(_06679_),
    .A2(_06680_),
    .B(_06681_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11723_ (.I(_06099_),
    .Z(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11724_ (.A1(_06675_),
    .A2(\register_file[8][16] ),
    .ZN(_06683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11725_ (.A1(_06682_),
    .A2(_06680_),
    .B(_06683_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11726_ (.I(_06103_),
    .Z(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11727_ (.A1(_06675_),
    .A2(\register_file[8][17] ),
    .ZN(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11728_ (.A1(_06684_),
    .A2(_06680_),
    .B(_06685_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11729_ (.I(_06107_),
    .Z(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11730_ (.I(_06639_),
    .Z(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11731_ (.A1(_06687_),
    .A2(\register_file[8][18] ),
    .ZN(_06688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11732_ (.A1(_06686_),
    .A2(_06680_),
    .B(_06688_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11733_ (.I(_06112_),
    .Z(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11734_ (.A1(_06687_),
    .A2(\register_file[8][19] ),
    .ZN(_06690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11735_ (.A1(_06689_),
    .A2(_06680_),
    .B(_06690_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11736_ (.I(_06116_),
    .Z(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11737_ (.I(_06655_),
    .Z(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11738_ (.A1(_06687_),
    .A2(\register_file[8][20] ),
    .ZN(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11739_ (.A1(_06691_),
    .A2(_06692_),
    .B(_06693_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11740_ (.I(_06121_),
    .Z(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11741_ (.A1(_06687_),
    .A2(\register_file[8][21] ),
    .ZN(_06695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11742_ (.A1(_06694_),
    .A2(_06692_),
    .B(_06695_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11743_ (.I(_06125_),
    .Z(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11744_ (.A1(_06687_),
    .A2(\register_file[8][22] ),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11745_ (.A1(_06696_),
    .A2(_06692_),
    .B(_06697_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11746_ (.I(_06129_),
    .Z(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11747_ (.I(_06639_),
    .Z(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11748_ (.A1(_06699_),
    .A2(\register_file[8][23] ),
    .ZN(_06700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11749_ (.A1(_06698_),
    .A2(_06692_),
    .B(_06700_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11750_ (.I(_06134_),
    .Z(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11751_ (.A1(_06699_),
    .A2(\register_file[8][24] ),
    .ZN(_06702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11752_ (.A1(_06701_),
    .A2(_06692_),
    .B(_06702_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11753_ (.I(_06138_),
    .Z(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11754_ (.I(_06655_),
    .Z(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11755_ (.A1(_06699_),
    .A2(\register_file[8][25] ),
    .ZN(_06705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11756_ (.A1(_06703_),
    .A2(_06704_),
    .B(_06705_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11757_ (.I(_06143_),
    .Z(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11758_ (.A1(_06699_),
    .A2(\register_file[8][26] ),
    .ZN(_06707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11759_ (.A1(_06706_),
    .A2(_06704_),
    .B(_06707_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11760_ (.I(_06147_),
    .Z(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11761_ (.A1(_06699_),
    .A2(\register_file[8][27] ),
    .ZN(_06709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11762_ (.A1(_06708_),
    .A2(_06704_),
    .B(_06709_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11763_ (.I(_06151_),
    .Z(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11764_ (.A1(_06640_),
    .A2(\register_file[8][28] ),
    .ZN(_06711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11765_ (.A1(_06710_),
    .A2(_06704_),
    .B(_06711_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11766_ (.I(_06155_),
    .Z(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11767_ (.A1(_06640_),
    .A2(\register_file[8][29] ),
    .ZN(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11768_ (.A1(_06712_),
    .A2(_06704_),
    .B(_06713_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11769_ (.I(_06159_),
    .Z(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11770_ (.A1(_06640_),
    .A2(\register_file[8][30] ),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11771_ (.A1(_06714_),
    .A2(_06643_),
    .B(_06715_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11772_ (.I(_06163_),
    .Z(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11773_ (.A1(_06640_),
    .A2(\register_file[8][31] ),
    .ZN(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11774_ (.A1(_06716_),
    .A2(_06643_),
    .B(_06717_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11775_ (.A1(_06266_),
    .A2(_03913_),
    .ZN(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11776_ (.I(_06718_),
    .Z(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11777_ (.I(_06719_),
    .Z(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11778_ (.I(_06718_),
    .Z(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11779_ (.I(_06721_),
    .Z(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11780_ (.A1(_06722_),
    .A2(\register_file[7][0] ),
    .ZN(_06723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11781_ (.A1(_06638_),
    .A2(_06720_),
    .B(_06723_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11782_ (.A1(_06722_),
    .A2(\register_file[7][1] ),
    .ZN(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11783_ (.A1(_06645_),
    .A2(_06720_),
    .B(_06724_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11784_ (.A1(_06722_),
    .A2(\register_file[7][2] ),
    .ZN(_06725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11785_ (.A1(_06647_),
    .A2(_06720_),
    .B(_06725_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11786_ (.I(_06721_),
    .Z(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11787_ (.A1(_06726_),
    .A2(\register_file[7][3] ),
    .ZN(_06727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11788_ (.A1(_06649_),
    .A2(_06720_),
    .B(_06727_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11789_ (.A1(_06726_),
    .A2(\register_file[7][4] ),
    .ZN(_06728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11790_ (.A1(_06652_),
    .A2(_06720_),
    .B(_06728_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11791_ (.I(_06721_),
    .Z(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11792_ (.I(_06729_),
    .Z(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11793_ (.A1(_06726_),
    .A2(\register_file[7][5] ),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11794_ (.A1(_06654_),
    .A2(_06730_),
    .B(_06731_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11795_ (.A1(_06726_),
    .A2(\register_file[7][6] ),
    .ZN(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11796_ (.A1(_06658_),
    .A2(_06730_),
    .B(_06732_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11797_ (.A1(_06726_),
    .A2(\register_file[7][7] ),
    .ZN(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11798_ (.A1(_06660_),
    .A2(_06730_),
    .B(_06733_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11799_ (.I(_06721_),
    .Z(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11800_ (.A1(_06734_),
    .A2(\register_file[7][8] ),
    .ZN(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11801_ (.A1(_06662_),
    .A2(_06730_),
    .B(_06735_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11802_ (.A1(_06734_),
    .A2(\register_file[7][9] ),
    .ZN(_06736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11803_ (.A1(_06665_),
    .A2(_06730_),
    .B(_06736_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11804_ (.I(_06729_),
    .Z(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11805_ (.A1(_06734_),
    .A2(\register_file[7][10] ),
    .ZN(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11806_ (.A1(_06667_),
    .A2(_06737_),
    .B(_06738_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11807_ (.A1(_06734_),
    .A2(\register_file[7][11] ),
    .ZN(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11808_ (.A1(_06670_),
    .A2(_06737_),
    .B(_06739_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11809_ (.A1(_06734_),
    .A2(\register_file[7][12] ),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11810_ (.A1(_06672_),
    .A2(_06737_),
    .B(_06740_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11811_ (.I(_06721_),
    .Z(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11812_ (.A1(_06741_),
    .A2(\register_file[7][13] ),
    .ZN(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11813_ (.A1(_06674_),
    .A2(_06737_),
    .B(_06742_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11814_ (.A1(_06741_),
    .A2(\register_file[7][14] ),
    .ZN(_06743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11815_ (.A1(_06677_),
    .A2(_06737_),
    .B(_06743_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11816_ (.I(_06729_),
    .Z(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11817_ (.A1(_06741_),
    .A2(\register_file[7][15] ),
    .ZN(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11818_ (.A1(_06679_),
    .A2(_06744_),
    .B(_06745_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11819_ (.A1(_06741_),
    .A2(\register_file[7][16] ),
    .ZN(_06746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11820_ (.A1(_06682_),
    .A2(_06744_),
    .B(_06746_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11821_ (.A1(_06741_),
    .A2(\register_file[7][17] ),
    .ZN(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11822_ (.A1(_06684_),
    .A2(_06744_),
    .B(_06747_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11823_ (.I(_06718_),
    .Z(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11824_ (.A1(_06748_),
    .A2(\register_file[7][18] ),
    .ZN(_06749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11825_ (.A1(_06686_),
    .A2(_06744_),
    .B(_06749_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11826_ (.A1(_06748_),
    .A2(\register_file[7][19] ),
    .ZN(_06750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11827_ (.A1(_06689_),
    .A2(_06744_),
    .B(_06750_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11828_ (.I(_06729_),
    .Z(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11829_ (.A1(_06748_),
    .A2(\register_file[7][20] ),
    .ZN(_06752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11830_ (.A1(_06691_),
    .A2(_06751_),
    .B(_06752_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11831_ (.A1(_06748_),
    .A2(\register_file[7][21] ),
    .ZN(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11832_ (.A1(_06694_),
    .A2(_06751_),
    .B(_06753_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11833_ (.A1(_06748_),
    .A2(\register_file[7][22] ),
    .ZN(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11834_ (.A1(_06696_),
    .A2(_06751_),
    .B(_06754_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11835_ (.I(_06718_),
    .Z(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11836_ (.A1(_06755_),
    .A2(\register_file[7][23] ),
    .ZN(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11837_ (.A1(_06698_),
    .A2(_06751_),
    .B(_06756_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11838_ (.A1(_06755_),
    .A2(\register_file[7][24] ),
    .ZN(_06757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11839_ (.A1(_06701_),
    .A2(_06751_),
    .B(_06757_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11840_ (.I(_06729_),
    .Z(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11841_ (.A1(_06755_),
    .A2(\register_file[7][25] ),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11842_ (.A1(_06703_),
    .A2(_06758_),
    .B(_06759_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11843_ (.A1(_06755_),
    .A2(\register_file[7][26] ),
    .ZN(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11844_ (.A1(_06706_),
    .A2(_06758_),
    .B(_06760_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11845_ (.A1(_06755_),
    .A2(\register_file[7][27] ),
    .ZN(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11846_ (.A1(_06708_),
    .A2(_06758_),
    .B(_06761_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11847_ (.A1(_06719_),
    .A2(\register_file[7][28] ),
    .ZN(_06762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11848_ (.A1(_06710_),
    .A2(_06758_),
    .B(_06762_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11849_ (.A1(_06719_),
    .A2(\register_file[7][29] ),
    .ZN(_06763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11850_ (.A1(_06712_),
    .A2(_06758_),
    .B(_06763_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11851_ (.A1(_06719_),
    .A2(\register_file[7][30] ),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11852_ (.A1(_06714_),
    .A2(_06722_),
    .B(_06764_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11853_ (.A1(_06719_),
    .A2(\register_file[7][31] ),
    .ZN(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11854_ (.A1(_06716_),
    .A2(_06722_),
    .B(_06765_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11855_ (.A1(_06024_),
    .A2(_03913_),
    .ZN(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11856_ (.I(_06766_),
    .Z(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11857_ (.I(_06767_),
    .Z(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11858_ (.I(_06766_),
    .Z(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11859_ (.I(_06769_),
    .Z(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11860_ (.A1(_06770_),
    .A2(\register_file[6][0] ),
    .ZN(_06771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11861_ (.A1(_06638_),
    .A2(_06768_),
    .B(_06771_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11862_ (.A1(_06770_),
    .A2(\register_file[6][1] ),
    .ZN(_06772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11863_ (.A1(_06645_),
    .A2(_06768_),
    .B(_06772_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11864_ (.A1(_06770_),
    .A2(\register_file[6][2] ),
    .ZN(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11865_ (.A1(_06647_),
    .A2(_06768_),
    .B(_06773_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11866_ (.I(_06769_),
    .Z(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11867_ (.A1(_06774_),
    .A2(\register_file[6][3] ),
    .ZN(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11868_ (.A1(_06649_),
    .A2(_06768_),
    .B(_06775_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11869_ (.A1(_06774_),
    .A2(\register_file[6][4] ),
    .ZN(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11870_ (.A1(_06652_),
    .A2(_06768_),
    .B(_06776_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11871_ (.I(_06769_),
    .Z(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11872_ (.I(_06777_),
    .Z(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11873_ (.A1(_06774_),
    .A2(\register_file[6][5] ),
    .ZN(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11874_ (.A1(_06654_),
    .A2(_06778_),
    .B(_06779_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11875_ (.A1(_06774_),
    .A2(\register_file[6][6] ),
    .ZN(_06780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11876_ (.A1(_06658_),
    .A2(_06778_),
    .B(_06780_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11877_ (.A1(_06774_),
    .A2(\register_file[6][7] ),
    .ZN(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11878_ (.A1(_06660_),
    .A2(_06778_),
    .B(_06781_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11879_ (.I(_06769_),
    .Z(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11880_ (.A1(_06782_),
    .A2(\register_file[6][8] ),
    .ZN(_06783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11881_ (.A1(_06662_),
    .A2(_06778_),
    .B(_06783_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11882_ (.A1(_06782_),
    .A2(\register_file[6][9] ),
    .ZN(_06784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11883_ (.A1(_06665_),
    .A2(_06778_),
    .B(_06784_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11884_ (.I(_06777_),
    .Z(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11885_ (.A1(_06782_),
    .A2(\register_file[6][10] ),
    .ZN(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11886_ (.A1(_06667_),
    .A2(_06785_),
    .B(_06786_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11887_ (.A1(_06782_),
    .A2(\register_file[6][11] ),
    .ZN(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11888_ (.A1(_06670_),
    .A2(_06785_),
    .B(_06787_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11889_ (.A1(_06782_),
    .A2(\register_file[6][12] ),
    .ZN(_06788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11890_ (.A1(_06672_),
    .A2(_06785_),
    .B(_06788_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11891_ (.I(_06769_),
    .Z(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11892_ (.A1(_06789_),
    .A2(\register_file[6][13] ),
    .ZN(_06790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11893_ (.A1(_06674_),
    .A2(_06785_),
    .B(_06790_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11894_ (.A1(_06789_),
    .A2(\register_file[6][14] ),
    .ZN(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11895_ (.A1(_06677_),
    .A2(_06785_),
    .B(_06791_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11896_ (.I(_06777_),
    .Z(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11897_ (.A1(_06789_),
    .A2(\register_file[6][15] ),
    .ZN(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11898_ (.A1(_06679_),
    .A2(_06792_),
    .B(_06793_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11899_ (.A1(_06789_),
    .A2(\register_file[6][16] ),
    .ZN(_06794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11900_ (.A1(_06682_),
    .A2(_06792_),
    .B(_06794_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11901_ (.A1(_06789_),
    .A2(\register_file[6][17] ),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11902_ (.A1(_06684_),
    .A2(_06792_),
    .B(_06795_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11903_ (.I(_06766_),
    .Z(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11904_ (.A1(_06796_),
    .A2(\register_file[6][18] ),
    .ZN(_06797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11905_ (.A1(_06686_),
    .A2(_06792_),
    .B(_06797_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11906_ (.A1(_06796_),
    .A2(\register_file[6][19] ),
    .ZN(_06798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11907_ (.A1(_06689_),
    .A2(_06792_),
    .B(_06798_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11908_ (.I(_06777_),
    .Z(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11909_ (.A1(_06796_),
    .A2(\register_file[6][20] ),
    .ZN(_06800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11910_ (.A1(_06691_),
    .A2(_06799_),
    .B(_06800_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11911_ (.A1(_06796_),
    .A2(\register_file[6][21] ),
    .ZN(_06801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11912_ (.A1(_06694_),
    .A2(_06799_),
    .B(_06801_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11913_ (.A1(_06796_),
    .A2(\register_file[6][22] ),
    .ZN(_06802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11914_ (.A1(_06696_),
    .A2(_06799_),
    .B(_06802_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11915_ (.I(_06766_),
    .Z(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11916_ (.A1(_06803_),
    .A2(\register_file[6][23] ),
    .ZN(_06804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11917_ (.A1(_06698_),
    .A2(_06799_),
    .B(_06804_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11918_ (.A1(_06803_),
    .A2(\register_file[6][24] ),
    .ZN(_06805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11919_ (.A1(_06701_),
    .A2(_06799_),
    .B(_06805_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11920_ (.I(_06777_),
    .Z(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11921_ (.A1(_06803_),
    .A2(\register_file[6][25] ),
    .ZN(_06807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11922_ (.A1(_06703_),
    .A2(_06806_),
    .B(_06807_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11923_ (.A1(_06803_),
    .A2(\register_file[6][26] ),
    .ZN(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11924_ (.A1(_06706_),
    .A2(_06806_),
    .B(_06808_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11925_ (.A1(_06803_),
    .A2(\register_file[6][27] ),
    .ZN(_06809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11926_ (.A1(_06708_),
    .A2(_06806_),
    .B(_06809_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11927_ (.A1(_06767_),
    .A2(\register_file[6][28] ),
    .ZN(_06810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11928_ (.A1(_06710_),
    .A2(_06806_),
    .B(_06810_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11929_ (.A1(_06767_),
    .A2(\register_file[6][29] ),
    .ZN(_06811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11930_ (.A1(_06712_),
    .A2(_06806_),
    .B(_06811_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11931_ (.A1(_06767_),
    .A2(\register_file[6][30] ),
    .ZN(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11932_ (.A1(_06714_),
    .A2(_06770_),
    .B(_06812_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11933_ (.A1(_06767_),
    .A2(\register_file[6][31] ),
    .ZN(_06813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11934_ (.A1(_06716_),
    .A2(_06770_),
    .B(_06813_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11935_ (.A1(_06317_),
    .A2(_03912_),
    .ZN(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11936_ (.I(_06814_),
    .Z(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11937_ (.I(_06815_),
    .Z(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11938_ (.I(_06814_),
    .Z(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11939_ (.I(_06817_),
    .Z(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11940_ (.A1(_06818_),
    .A2(\register_file[5][0] ),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11941_ (.A1(_06638_),
    .A2(_06816_),
    .B(_06819_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11942_ (.A1(_06818_),
    .A2(\register_file[5][1] ),
    .ZN(_06820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11943_ (.A1(_06645_),
    .A2(_06816_),
    .B(_06820_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11944_ (.A1(_06818_),
    .A2(\register_file[5][2] ),
    .ZN(_06821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11945_ (.A1(_06647_),
    .A2(_06816_),
    .B(_06821_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11946_ (.I(_06817_),
    .Z(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11947_ (.A1(_06822_),
    .A2(\register_file[5][3] ),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11948_ (.A1(_06649_),
    .A2(_06816_),
    .B(_06823_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11949_ (.A1(_06822_),
    .A2(\register_file[5][4] ),
    .ZN(_06824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11950_ (.A1(_06652_),
    .A2(_06816_),
    .B(_06824_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11951_ (.I(_06817_),
    .Z(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11952_ (.I(_06825_),
    .Z(_06826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11953_ (.A1(_06822_),
    .A2(\register_file[5][5] ),
    .ZN(_06827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11954_ (.A1(_06654_),
    .A2(_06826_),
    .B(_06827_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11955_ (.A1(_06822_),
    .A2(\register_file[5][6] ),
    .ZN(_06828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11956_ (.A1(_06658_),
    .A2(_06826_),
    .B(_06828_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11957_ (.A1(_06822_),
    .A2(\register_file[5][7] ),
    .ZN(_06829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11958_ (.A1(_06660_),
    .A2(_06826_),
    .B(_06829_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11959_ (.I(_06817_),
    .Z(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11960_ (.A1(_06830_),
    .A2(\register_file[5][8] ),
    .ZN(_06831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11961_ (.A1(_06662_),
    .A2(_06826_),
    .B(_06831_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11962_ (.A1(_06830_),
    .A2(\register_file[5][9] ),
    .ZN(_06832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11963_ (.A1(_06665_),
    .A2(_06826_),
    .B(_06832_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11964_ (.I(_06825_),
    .Z(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11965_ (.A1(_06830_),
    .A2(\register_file[5][10] ),
    .ZN(_06834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11966_ (.A1(_06667_),
    .A2(_06833_),
    .B(_06834_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11967_ (.A1(_06830_),
    .A2(\register_file[5][11] ),
    .ZN(_06835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11968_ (.A1(_06670_),
    .A2(_06833_),
    .B(_06835_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11969_ (.A1(_06830_),
    .A2(\register_file[5][12] ),
    .ZN(_06836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11970_ (.A1(_06672_),
    .A2(_06833_),
    .B(_06836_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11971_ (.I(_06817_),
    .Z(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11972_ (.A1(_06837_),
    .A2(\register_file[5][13] ),
    .ZN(_06838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11973_ (.A1(_06674_),
    .A2(_06833_),
    .B(_06838_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11974_ (.A1(_06837_),
    .A2(\register_file[5][14] ),
    .ZN(_06839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11975_ (.A1(_06677_),
    .A2(_06833_),
    .B(_06839_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11976_ (.I(_06825_),
    .Z(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11977_ (.A1(_06837_),
    .A2(\register_file[5][15] ),
    .ZN(_06841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11978_ (.A1(_06679_),
    .A2(_06840_),
    .B(_06841_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11979_ (.A1(_06837_),
    .A2(\register_file[5][16] ),
    .ZN(_06842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11980_ (.A1(_06682_),
    .A2(_06840_),
    .B(_06842_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11981_ (.A1(_06837_),
    .A2(\register_file[5][17] ),
    .ZN(_06843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11982_ (.A1(_06684_),
    .A2(_06840_),
    .B(_06843_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11983_ (.I(_06814_),
    .Z(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11984_ (.A1(_06844_),
    .A2(\register_file[5][18] ),
    .ZN(_06845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11985_ (.A1(_06686_),
    .A2(_06840_),
    .B(_06845_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11986_ (.A1(_06844_),
    .A2(\register_file[5][19] ),
    .ZN(_06846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11987_ (.A1(_06689_),
    .A2(_06840_),
    .B(_06846_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11988_ (.I(_06825_),
    .Z(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11989_ (.A1(_06844_),
    .A2(\register_file[5][20] ),
    .ZN(_06848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11990_ (.A1(_06691_),
    .A2(_06847_),
    .B(_06848_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11991_ (.A1(_06844_),
    .A2(\register_file[5][21] ),
    .ZN(_06849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11992_ (.A1(_06694_),
    .A2(_06847_),
    .B(_06849_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11993_ (.A1(_06844_),
    .A2(\register_file[5][22] ),
    .ZN(_06850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11994_ (.A1(_06696_),
    .A2(_06847_),
    .B(_06850_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11995_ (.I(_06814_),
    .Z(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11996_ (.A1(_06851_),
    .A2(\register_file[5][23] ),
    .ZN(_06852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11997_ (.A1(_06698_),
    .A2(_06847_),
    .B(_06852_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11998_ (.A1(_06851_),
    .A2(\register_file[5][24] ),
    .ZN(_06853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11999_ (.A1(_06701_),
    .A2(_06847_),
    .B(_06853_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12000_ (.I(_06825_),
    .Z(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12001_ (.A1(_06851_),
    .A2(\register_file[5][25] ),
    .ZN(_06855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12002_ (.A1(_06703_),
    .A2(_06854_),
    .B(_06855_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12003_ (.A1(_06851_),
    .A2(\register_file[5][26] ),
    .ZN(_06856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12004_ (.A1(_06706_),
    .A2(_06854_),
    .B(_06856_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12005_ (.A1(_06851_),
    .A2(\register_file[5][27] ),
    .ZN(_06857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12006_ (.A1(_06708_),
    .A2(_06854_),
    .B(_06857_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12007_ (.A1(_06815_),
    .A2(\register_file[5][28] ),
    .ZN(_06858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12008_ (.A1(_06710_),
    .A2(_06854_),
    .B(_06858_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12009_ (.A1(_06815_),
    .A2(\register_file[5][29] ),
    .ZN(_06859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12010_ (.A1(_06712_),
    .A2(_06854_),
    .B(_06859_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12011_ (.A1(_06815_),
    .A2(\register_file[5][30] ),
    .ZN(_06860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12012_ (.A1(_06714_),
    .A2(_06818_),
    .B(_06860_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12013_ (.A1(_06815_),
    .A2(\register_file[5][31] ),
    .ZN(_06861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12014_ (.A1(_06716_),
    .A2(_06818_),
    .B(_06861_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12015_ (.A1(_03911_),
    .A2(_06214_),
    .ZN(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12016_ (.I(_06862_),
    .Z(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12017_ (.I(_06863_),
    .Z(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12018_ (.I(_06862_),
    .Z(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12019_ (.I(_06865_),
    .Z(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12020_ (.A1(_06866_),
    .A2(net11),
    .ZN(_06867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12021_ (.A1(_01163_),
    .A2(_06864_),
    .B(_06867_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12022_ (.A1(_06866_),
    .A2(net22),
    .ZN(_06868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12023_ (.A1(_01268_),
    .A2(_06864_),
    .B(_06868_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12024_ (.A1(_06866_),
    .A2(net33),
    .ZN(_06869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12025_ (.A1(_01358_),
    .A2(_06864_),
    .B(_06869_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12026_ (.I(_06865_),
    .Z(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12027_ (.A1(_06870_),
    .A2(net36),
    .ZN(_06871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12028_ (.A1(_01446_),
    .A2(_06864_),
    .B(_06871_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12029_ (.A1(_06870_),
    .A2(net37),
    .ZN(_06872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12030_ (.A1(_01532_),
    .A2(_06864_),
    .B(_06872_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12031_ (.I(_06865_),
    .Z(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12032_ (.I(_06873_),
    .Z(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12033_ (.A1(_06870_),
    .A2(net38),
    .ZN(_06875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12034_ (.A1(_01616_),
    .A2(_06874_),
    .B(_06875_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12035_ (.A1(_06870_),
    .A2(net39),
    .ZN(_06876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12036_ (.A1(_01704_),
    .A2(_06874_),
    .B(_06876_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12037_ (.A1(_06870_),
    .A2(net40),
    .ZN(_06877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12038_ (.A1(_01789_),
    .A2(_06874_),
    .B(_06877_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12039_ (.I(_06865_),
    .Z(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12040_ (.A1(_06878_),
    .A2(net41),
    .ZN(_06879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12041_ (.A1(_01874_),
    .A2(_06874_),
    .B(_06879_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12042_ (.A1(_06878_),
    .A2(net42),
    .ZN(_06880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12043_ (.A1(_01955_),
    .A2(_06874_),
    .B(_06880_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12044_ (.I(_06873_),
    .Z(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12045_ (.A1(_06878_),
    .A2(net12),
    .ZN(_06882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12046_ (.A1(_02038_),
    .A2(_06881_),
    .B(_06882_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12047_ (.A1(_06878_),
    .A2(net13),
    .ZN(_06883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12048_ (.A1(_02122_),
    .A2(_06881_),
    .B(_06883_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12049_ (.A1(_06878_),
    .A2(net14),
    .ZN(_06884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12050_ (.A1(_02206_),
    .A2(_06881_),
    .B(_06884_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12051_ (.I(_06865_),
    .Z(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12052_ (.A1(_06885_),
    .A2(net15),
    .ZN(_06886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12053_ (.A1(_02291_),
    .A2(_06881_),
    .B(_06886_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12054_ (.A1(_06885_),
    .A2(net16),
    .ZN(_06887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12055_ (.A1(_02372_),
    .A2(_06881_),
    .B(_06887_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12056_ (.I(_06873_),
    .Z(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12057_ (.A1(_06885_),
    .A2(net17),
    .ZN(_06889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12058_ (.A1(_02455_),
    .A2(_06888_),
    .B(_06889_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12059_ (.A1(_06885_),
    .A2(net18),
    .ZN(_06890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12060_ (.A1(_02539_),
    .A2(_06888_),
    .B(_06890_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12061_ (.A1(_06885_),
    .A2(net19),
    .ZN(_06891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12062_ (.A1(_02623_),
    .A2(_06888_),
    .B(_06891_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12063_ (.I(_06862_),
    .Z(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12064_ (.A1(_06892_),
    .A2(net20),
    .ZN(_06893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12065_ (.A1(_02706_),
    .A2(_06888_),
    .B(_06893_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12066_ (.A1(_06892_),
    .A2(net21),
    .ZN(_06894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12067_ (.A1(_02787_),
    .A2(_06888_),
    .B(_06894_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12068_ (.I(_06873_),
    .Z(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12069_ (.A1(_06892_),
    .A2(net23),
    .ZN(_06896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12070_ (.A1(_02870_),
    .A2(_06895_),
    .B(_06896_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12071_ (.A1(_06892_),
    .A2(net24),
    .ZN(_06897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12072_ (.A1(_02955_),
    .A2(_06895_),
    .B(_06897_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12073_ (.A1(_06892_),
    .A2(net25),
    .ZN(_06898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12074_ (.A1(_03040_),
    .A2(_06895_),
    .B(_06898_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12075_ (.I(_06862_),
    .Z(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12076_ (.A1(_06899_),
    .A2(net26),
    .ZN(_06900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12077_ (.A1(_03123_),
    .A2(_06895_),
    .B(_06900_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12078_ (.A1(_06899_),
    .A2(net27),
    .ZN(_06901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12079_ (.A1(_03204_),
    .A2(_06895_),
    .B(_06901_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12080_ (.I(_06873_),
    .Z(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12081_ (.A1(_06899_),
    .A2(net28),
    .ZN(_06903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12082_ (.A1(_03287_),
    .A2(_06902_),
    .B(_06903_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12083_ (.A1(_06899_),
    .A2(net29),
    .ZN(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12084_ (.A1(_03371_),
    .A2(_06902_),
    .B(_06904_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12085_ (.A1(_06899_),
    .A2(net30),
    .ZN(_06905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12086_ (.A1(_03448_),
    .A2(_06902_),
    .B(_06905_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12087_ (.A1(_06863_),
    .A2(net31),
    .ZN(_06906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12088_ (.A1(_03521_),
    .A2(_06902_),
    .B(_06906_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12089_ (.A1(_06863_),
    .A2(net32),
    .ZN(_06907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12090_ (.A1(_03593_),
    .A2(_06902_),
    .B(_06907_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12091_ (.A1(_06863_),
    .A2(net34),
    .ZN(_06908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12092_ (.A1(_03666_),
    .A2(_06866_),
    .B(_06908_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12093_ (.A1(_06863_),
    .A2(net35),
    .ZN(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12094_ (.A1(_03686_),
    .A2(_06866_),
    .B(_06909_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12095_ (.A1(_06266_),
    .A2(_03927_),
    .ZN(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12096_ (.I(_06910_),
    .Z(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12097_ (.I(_06911_),
    .Z(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12098_ (.I(_06910_),
    .Z(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12099_ (.I(_06913_),
    .Z(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12100_ (.A1(_06914_),
    .A2(\register_file[3][0] ),
    .ZN(_06915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12101_ (.A1(_06638_),
    .A2(_06912_),
    .B(_06915_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12102_ (.A1(_06914_),
    .A2(\register_file[3][1] ),
    .ZN(_06916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12103_ (.A1(_06645_),
    .A2(_06912_),
    .B(_06916_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12104_ (.A1(_06914_),
    .A2(\register_file[3][2] ),
    .ZN(_06917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12105_ (.A1(_06647_),
    .A2(_06912_),
    .B(_06917_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12106_ (.I(_06913_),
    .Z(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12107_ (.A1(_06918_),
    .A2(\register_file[3][3] ),
    .ZN(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12108_ (.A1(_06649_),
    .A2(_06912_),
    .B(_06919_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12109_ (.A1(_06918_),
    .A2(\register_file[3][4] ),
    .ZN(_06920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12110_ (.A1(_06652_),
    .A2(_06912_),
    .B(_06920_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12111_ (.I(_06913_),
    .Z(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12112_ (.I(_06921_),
    .Z(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12113_ (.A1(_06918_),
    .A2(\register_file[3][5] ),
    .ZN(_06923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12114_ (.A1(_06654_),
    .A2(_06922_),
    .B(_06923_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12115_ (.A1(_06918_),
    .A2(\register_file[3][6] ),
    .ZN(_06924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12116_ (.A1(_06658_),
    .A2(_06922_),
    .B(_06924_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12117_ (.A1(_06918_),
    .A2(\register_file[3][7] ),
    .ZN(_06925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12118_ (.A1(_06660_),
    .A2(_06922_),
    .B(_06925_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12119_ (.I(_06913_),
    .Z(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12120_ (.A1(_06926_),
    .A2(\register_file[3][8] ),
    .ZN(_06927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12121_ (.A1(_06662_),
    .A2(_06922_),
    .B(_06927_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12122_ (.A1(_06926_),
    .A2(\register_file[3][9] ),
    .ZN(_06928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12123_ (.A1(_06665_),
    .A2(_06922_),
    .B(_06928_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12124_ (.I(_06921_),
    .Z(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12125_ (.A1(_06926_),
    .A2(\register_file[3][10] ),
    .ZN(_06930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12126_ (.A1(_06667_),
    .A2(_06929_),
    .B(_06930_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12127_ (.A1(_06926_),
    .A2(\register_file[3][11] ),
    .ZN(_06931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12128_ (.A1(_06670_),
    .A2(_06929_),
    .B(_06931_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12129_ (.A1(_06926_),
    .A2(\register_file[3][12] ),
    .ZN(_06932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12130_ (.A1(_06672_),
    .A2(_06929_),
    .B(_06932_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12131_ (.I(_06913_),
    .Z(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12132_ (.A1(_06933_),
    .A2(\register_file[3][13] ),
    .ZN(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12133_ (.A1(_06674_),
    .A2(_06929_),
    .B(_06934_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12134_ (.A1(_06933_),
    .A2(\register_file[3][14] ),
    .ZN(_06935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12135_ (.A1(_06677_),
    .A2(_06929_),
    .B(_06935_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12136_ (.I(_06921_),
    .Z(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12137_ (.A1(_06933_),
    .A2(\register_file[3][15] ),
    .ZN(_06937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12138_ (.A1(_06679_),
    .A2(_06936_),
    .B(_06937_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12139_ (.A1(_06933_),
    .A2(\register_file[3][16] ),
    .ZN(_06938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12140_ (.A1(_06682_),
    .A2(_06936_),
    .B(_06938_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12141_ (.A1(_06933_),
    .A2(\register_file[3][17] ),
    .ZN(_06939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12142_ (.A1(_06684_),
    .A2(_06936_),
    .B(_06939_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12143_ (.I(_06910_),
    .Z(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12144_ (.A1(_06940_),
    .A2(\register_file[3][18] ),
    .ZN(_06941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12145_ (.A1(_06686_),
    .A2(_06936_),
    .B(_06941_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12146_ (.A1(_06940_),
    .A2(\register_file[3][19] ),
    .ZN(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12147_ (.A1(_06689_),
    .A2(_06936_),
    .B(_06942_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12148_ (.I(_06921_),
    .Z(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12149_ (.A1(_06940_),
    .A2(\register_file[3][20] ),
    .ZN(_06944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12150_ (.A1(_06691_),
    .A2(_06943_),
    .B(_06944_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12151_ (.A1(_06940_),
    .A2(\register_file[3][21] ),
    .ZN(_06945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12152_ (.A1(_06694_),
    .A2(_06943_),
    .B(_06945_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12153_ (.A1(_06940_),
    .A2(\register_file[3][22] ),
    .ZN(_06946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12154_ (.A1(_06696_),
    .A2(_06943_),
    .B(_06946_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12155_ (.I(_06910_),
    .Z(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12156_ (.A1(_06947_),
    .A2(\register_file[3][23] ),
    .ZN(_06948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12157_ (.A1(_06698_),
    .A2(_06943_),
    .B(_06948_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12158_ (.A1(_06947_),
    .A2(\register_file[3][24] ),
    .ZN(_06949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12159_ (.A1(_06701_),
    .A2(_06943_),
    .B(_06949_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12160_ (.I(_06921_),
    .Z(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12161_ (.A1(_06947_),
    .A2(\register_file[3][25] ),
    .ZN(_06951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12162_ (.A1(_06703_),
    .A2(_06950_),
    .B(_06951_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12163_ (.A1(_06947_),
    .A2(\register_file[3][26] ),
    .ZN(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12164_ (.A1(_06706_),
    .A2(_06950_),
    .B(_06952_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12165_ (.A1(_06947_),
    .A2(\register_file[3][27] ),
    .ZN(_06953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12166_ (.A1(_06708_),
    .A2(_06950_),
    .B(_06953_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12167_ (.A1(_06911_),
    .A2(\register_file[3][28] ),
    .ZN(_06954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12168_ (.A1(_06710_),
    .A2(_06950_),
    .B(_06954_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12169_ (.A1(_06911_),
    .A2(\register_file[3][29] ),
    .ZN(_06955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12170_ (.A1(_06712_),
    .A2(_06950_),
    .B(_06955_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12171_ (.A1(_06911_),
    .A2(\register_file[3][30] ),
    .ZN(_06956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12172_ (.A1(_06714_),
    .A2(_06914_),
    .B(_06956_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12173_ (.A1(_06911_),
    .A2(\register_file[3][31] ),
    .ZN(_06957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12174_ (.A1(_06716_),
    .A2(_06914_),
    .B(_06957_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12175_ (.I(_06020_),
    .Z(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12176_ (.A1(_06265_),
    .A2(_03815_),
    .ZN(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12177_ (.I(_06959_),
    .Z(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12178_ (.I(_06960_),
    .Z(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12179_ (.I(_06959_),
    .Z(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12180_ (.I(_06962_),
    .Z(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12181_ (.A1(_06963_),
    .A2(\register_file[31][0] ),
    .ZN(_06964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12182_ (.A1(_06958_),
    .A2(_06961_),
    .B(_06964_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12183_ (.I(_06032_),
    .Z(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12184_ (.A1(_06963_),
    .A2(\register_file[31][1] ),
    .ZN(_06966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12185_ (.A1(_06965_),
    .A2(_06961_),
    .B(_06966_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12186_ (.I(_06036_),
    .Z(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12187_ (.A1(_06963_),
    .A2(\register_file[31][2] ),
    .ZN(_06968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12188_ (.A1(_06967_),
    .A2(_06961_),
    .B(_06968_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12189_ (.I(_06040_),
    .Z(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12190_ (.I(_06962_),
    .Z(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12191_ (.A1(_06970_),
    .A2(\register_file[31][3] ),
    .ZN(_06971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12192_ (.A1(_06969_),
    .A2(_06961_),
    .B(_06971_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12193_ (.I(_06045_),
    .Z(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12194_ (.A1(_06970_),
    .A2(\register_file[31][4] ),
    .ZN(_06973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12195_ (.A1(_06972_),
    .A2(_06961_),
    .B(_06973_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12196_ (.I(_06049_),
    .Z(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12197_ (.I(_06962_),
    .Z(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12198_ (.I(_06975_),
    .Z(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12199_ (.A1(_06970_),
    .A2(\register_file[31][5] ),
    .ZN(_06977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12200_ (.A1(_06974_),
    .A2(_06976_),
    .B(_06977_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12201_ (.I(_06055_),
    .Z(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12202_ (.A1(_06970_),
    .A2(\register_file[31][6] ),
    .ZN(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12203_ (.A1(_06978_),
    .A2(_06976_),
    .B(_06979_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12204_ (.I(_06059_),
    .Z(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12205_ (.A1(_06970_),
    .A2(\register_file[31][7] ),
    .ZN(_06981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12206_ (.A1(_06980_),
    .A2(_06976_),
    .B(_06981_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12207_ (.I(_06063_),
    .Z(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12208_ (.I(_06962_),
    .Z(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12209_ (.A1(_06983_),
    .A2(\register_file[31][8] ),
    .ZN(_06984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12210_ (.A1(_06982_),
    .A2(_06976_),
    .B(_06984_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12211_ (.I(_06068_),
    .Z(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12212_ (.A1(_06983_),
    .A2(\register_file[31][9] ),
    .ZN(_06986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12213_ (.A1(_06985_),
    .A2(_06976_),
    .B(_06986_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12214_ (.I(_06072_),
    .Z(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12215_ (.I(_06975_),
    .Z(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12216_ (.A1(_06983_),
    .A2(\register_file[31][10] ),
    .ZN(_06989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12217_ (.A1(_06987_),
    .A2(_06988_),
    .B(_06989_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12218_ (.I(_06077_),
    .Z(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12219_ (.A1(_06983_),
    .A2(\register_file[31][11] ),
    .ZN(_06991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12220_ (.A1(_06990_),
    .A2(_06988_),
    .B(_06991_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12221_ (.I(_06081_),
    .Z(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12222_ (.A1(_06983_),
    .A2(\register_file[31][12] ),
    .ZN(_06993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12223_ (.A1(_06992_),
    .A2(_06988_),
    .B(_06993_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12224_ (.I(_06085_),
    .Z(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12225_ (.I(_06962_),
    .Z(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12226_ (.A1(_06995_),
    .A2(\register_file[31][13] ),
    .ZN(_06996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12227_ (.A1(_06994_),
    .A2(_06988_),
    .B(_06996_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12228_ (.I(_06090_),
    .Z(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12229_ (.A1(_06995_),
    .A2(\register_file[31][14] ),
    .ZN(_06998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12230_ (.A1(_06997_),
    .A2(_06988_),
    .B(_06998_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12231_ (.I(_06094_),
    .Z(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12232_ (.I(_06975_),
    .Z(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12233_ (.A1(_06995_),
    .A2(\register_file[31][15] ),
    .ZN(_07001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12234_ (.A1(_06999_),
    .A2(_07000_),
    .B(_07001_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12235_ (.I(_06099_),
    .Z(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12236_ (.A1(_06995_),
    .A2(\register_file[31][16] ),
    .ZN(_07003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12237_ (.A1(_07002_),
    .A2(_07000_),
    .B(_07003_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12238_ (.I(_06103_),
    .Z(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12239_ (.A1(_06995_),
    .A2(\register_file[31][17] ),
    .ZN(_07005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12240_ (.A1(_07004_),
    .A2(_07000_),
    .B(_07005_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12241_ (.I(_06107_),
    .Z(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12242_ (.I(_06959_),
    .Z(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12243_ (.A1(_07007_),
    .A2(\register_file[31][18] ),
    .ZN(_07008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12244_ (.A1(_07006_),
    .A2(_07000_),
    .B(_07008_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12245_ (.I(_06112_),
    .Z(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12246_ (.A1(_07007_),
    .A2(\register_file[31][19] ),
    .ZN(_07010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12247_ (.A1(_07009_),
    .A2(_07000_),
    .B(_07010_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12248_ (.I(_06116_),
    .Z(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12249_ (.I(_06975_),
    .Z(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12250_ (.A1(_07007_),
    .A2(\register_file[31][20] ),
    .ZN(_07013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12251_ (.A1(_07011_),
    .A2(_07012_),
    .B(_07013_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12252_ (.I(_06121_),
    .Z(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12253_ (.A1(_07007_),
    .A2(\register_file[31][21] ),
    .ZN(_07015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12254_ (.A1(_07014_),
    .A2(_07012_),
    .B(_07015_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12255_ (.I(_06125_),
    .Z(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12256_ (.A1(_07007_),
    .A2(\register_file[31][22] ),
    .ZN(_07017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12257_ (.A1(_07016_),
    .A2(_07012_),
    .B(_07017_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12258_ (.I(_06129_),
    .Z(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12259_ (.I(_06959_),
    .Z(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12260_ (.A1(_07019_),
    .A2(\register_file[31][23] ),
    .ZN(_07020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12261_ (.A1(_07018_),
    .A2(_07012_),
    .B(_07020_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12262_ (.I(_06134_),
    .Z(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12263_ (.A1(_07019_),
    .A2(\register_file[31][24] ),
    .ZN(_07022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12264_ (.A1(_07021_),
    .A2(_07012_),
    .B(_07022_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12265_ (.I(_06138_),
    .Z(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12266_ (.I(_06975_),
    .Z(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12267_ (.A1(_07019_),
    .A2(\register_file[31][25] ),
    .ZN(_07025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12268_ (.A1(_07023_),
    .A2(_07024_),
    .B(_07025_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12269_ (.I(_06143_),
    .Z(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12270_ (.A1(_07019_),
    .A2(\register_file[31][26] ),
    .ZN(_07027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12271_ (.A1(_07026_),
    .A2(_07024_),
    .B(_07027_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12272_ (.I(_06147_),
    .Z(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12273_ (.A1(_07019_),
    .A2(\register_file[31][27] ),
    .ZN(_07029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12274_ (.A1(_07028_),
    .A2(_07024_),
    .B(_07029_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12275_ (.I(_06151_),
    .Z(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12276_ (.A1(_06960_),
    .A2(\register_file[31][28] ),
    .ZN(_07031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12277_ (.A1(_07030_),
    .A2(_07024_),
    .B(_07031_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12278_ (.I(_06155_),
    .Z(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12279_ (.A1(_06960_),
    .A2(\register_file[31][29] ),
    .ZN(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12280_ (.A1(_07032_),
    .A2(_07024_),
    .B(_07033_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12281_ (.I(_06159_),
    .Z(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12282_ (.A1(_06960_),
    .A2(\register_file[31][30] ),
    .ZN(_07035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12283_ (.A1(_07034_),
    .A2(_06963_),
    .B(_07035_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12284_ (.I(_06163_),
    .Z(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12285_ (.A1(_06960_),
    .A2(\register_file[31][31] ),
    .ZN(_07037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12286_ (.A1(_07036_),
    .A2(_06963_),
    .B(_07037_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12287_ (.A1(_06317_),
    .A2(_03794_),
    .ZN(_07038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12288_ (.I(_07038_),
    .Z(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12289_ (.I(_07039_),
    .Z(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12290_ (.I(_07038_),
    .Z(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12291_ (.I(_07041_),
    .Z(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12292_ (.A1(_07042_),
    .A2(\register_file[25][0] ),
    .ZN(_07043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12293_ (.A1(_06958_),
    .A2(_07040_),
    .B(_07043_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12294_ (.A1(_07042_),
    .A2(\register_file[25][1] ),
    .ZN(_07044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12295_ (.A1(_06965_),
    .A2(_07040_),
    .B(_07044_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12296_ (.A1(_07042_),
    .A2(\register_file[25][2] ),
    .ZN(_07045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12297_ (.A1(_06967_),
    .A2(_07040_),
    .B(_07045_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12298_ (.I(_07041_),
    .Z(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12299_ (.A1(_07046_),
    .A2(\register_file[25][3] ),
    .ZN(_07047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12300_ (.A1(_06969_),
    .A2(_07040_),
    .B(_07047_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12301_ (.A1(_07046_),
    .A2(\register_file[25][4] ),
    .ZN(_07048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12302_ (.A1(_06972_),
    .A2(_07040_),
    .B(_07048_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12303_ (.I(_07041_),
    .Z(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12304_ (.I(_07049_),
    .Z(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12305_ (.A1(_07046_),
    .A2(\register_file[25][5] ),
    .ZN(_07051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12306_ (.A1(_06974_),
    .A2(_07050_),
    .B(_07051_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12307_ (.A1(_07046_),
    .A2(\register_file[25][6] ),
    .ZN(_07052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12308_ (.A1(_06978_),
    .A2(_07050_),
    .B(_07052_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12309_ (.A1(_07046_),
    .A2(\register_file[25][7] ),
    .ZN(_07053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12310_ (.A1(_06980_),
    .A2(_07050_),
    .B(_07053_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12311_ (.I(_07041_),
    .Z(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12312_ (.A1(_07054_),
    .A2(\register_file[25][8] ),
    .ZN(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12313_ (.A1(_06982_),
    .A2(_07050_),
    .B(_07055_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12314_ (.A1(_07054_),
    .A2(\register_file[25][9] ),
    .ZN(_07056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12315_ (.A1(_06985_),
    .A2(_07050_),
    .B(_07056_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12316_ (.I(_07049_),
    .Z(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12317_ (.A1(_07054_),
    .A2(\register_file[25][10] ),
    .ZN(_07058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12318_ (.A1(_06987_),
    .A2(_07057_),
    .B(_07058_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12319_ (.A1(_07054_),
    .A2(\register_file[25][11] ),
    .ZN(_07059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12320_ (.A1(_06990_),
    .A2(_07057_),
    .B(_07059_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12321_ (.A1(_07054_),
    .A2(\register_file[25][12] ),
    .ZN(_07060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12322_ (.A1(_06992_),
    .A2(_07057_),
    .B(_07060_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12323_ (.I(_07041_),
    .Z(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12324_ (.A1(_07061_),
    .A2(\register_file[25][13] ),
    .ZN(_07062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12325_ (.A1(_06994_),
    .A2(_07057_),
    .B(_07062_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12326_ (.A1(_07061_),
    .A2(\register_file[25][14] ),
    .ZN(_07063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12327_ (.A1(_06997_),
    .A2(_07057_),
    .B(_07063_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12328_ (.I(_07049_),
    .Z(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12329_ (.A1(_07061_),
    .A2(\register_file[25][15] ),
    .ZN(_07065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12330_ (.A1(_06999_),
    .A2(_07064_),
    .B(_07065_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12331_ (.A1(_07061_),
    .A2(\register_file[25][16] ),
    .ZN(_07066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12332_ (.A1(_07002_),
    .A2(_07064_),
    .B(_07066_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12333_ (.A1(_07061_),
    .A2(\register_file[25][17] ),
    .ZN(_07067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12334_ (.A1(_07004_),
    .A2(_07064_),
    .B(_07067_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12335_ (.I(_07038_),
    .Z(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12336_ (.A1(_07068_),
    .A2(\register_file[25][18] ),
    .ZN(_07069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12337_ (.A1(_07006_),
    .A2(_07064_),
    .B(_07069_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12338_ (.A1(_07068_),
    .A2(\register_file[25][19] ),
    .ZN(_07070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12339_ (.A1(_07009_),
    .A2(_07064_),
    .B(_07070_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12340_ (.I(_07049_),
    .Z(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12341_ (.A1(_07068_),
    .A2(\register_file[25][20] ),
    .ZN(_07072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12342_ (.A1(_07011_),
    .A2(_07071_),
    .B(_07072_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12343_ (.A1(_07068_),
    .A2(\register_file[25][21] ),
    .ZN(_07073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12344_ (.A1(_07014_),
    .A2(_07071_),
    .B(_07073_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12345_ (.A1(_07068_),
    .A2(\register_file[25][22] ),
    .ZN(_07074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12346_ (.A1(_07016_),
    .A2(_07071_),
    .B(_07074_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12347_ (.I(_07038_),
    .Z(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12348_ (.A1(_07075_),
    .A2(\register_file[25][23] ),
    .ZN(_07076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12349_ (.A1(_07018_),
    .A2(_07071_),
    .B(_07076_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12350_ (.A1(_07075_),
    .A2(\register_file[25][24] ),
    .ZN(_07077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12351_ (.A1(_07021_),
    .A2(_07071_),
    .B(_07077_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12352_ (.I(_07049_),
    .Z(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12353_ (.A1(_07075_),
    .A2(\register_file[25][25] ),
    .ZN(_07079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12354_ (.A1(_07023_),
    .A2(_07078_),
    .B(_07079_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12355_ (.A1(_07075_),
    .A2(\register_file[25][26] ),
    .ZN(_07080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12356_ (.A1(_07026_),
    .A2(_07078_),
    .B(_07080_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12357_ (.A1(_07075_),
    .A2(\register_file[25][27] ),
    .ZN(_07081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12358_ (.A1(_07028_),
    .A2(_07078_),
    .B(_07081_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12359_ (.A1(_07039_),
    .A2(\register_file[25][28] ),
    .ZN(_07082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12360_ (.A1(_07030_),
    .A2(_07078_),
    .B(_07082_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12361_ (.A1(_07039_),
    .A2(\register_file[25][29] ),
    .ZN(_07083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12362_ (.A1(_07032_),
    .A2(_07078_),
    .B(_07083_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12363_ (.A1(_07039_),
    .A2(\register_file[25][30] ),
    .ZN(_07084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12364_ (.A1(_07034_),
    .A2(_07042_),
    .B(_07084_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12365_ (.A1(_07039_),
    .A2(\register_file[25][31] ),
    .ZN(_07085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12366_ (.A1(_07036_),
    .A2(_07042_),
    .B(_07085_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12367_ (.A1(_04067_),
    .A2(_06215_),
    .ZN(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12368_ (.I(_07086_),
    .Z(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12369_ (.I(_07087_),
    .Z(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12370_ (.I(_07086_),
    .Z(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12371_ (.I(_07089_),
    .Z(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12372_ (.A1(_07090_),
    .A2(\register_file[24][0] ),
    .ZN(_07091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12373_ (.A1(_06958_),
    .A2(_07088_),
    .B(_07091_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12374_ (.A1(_07090_),
    .A2(\register_file[24][1] ),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12375_ (.A1(_06965_),
    .A2(_07088_),
    .B(_07092_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12376_ (.A1(_07090_),
    .A2(\register_file[24][2] ),
    .ZN(_07093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12377_ (.A1(_06967_),
    .A2(_07088_),
    .B(_07093_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12378_ (.I(_07089_),
    .Z(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12379_ (.A1(_07094_),
    .A2(\register_file[24][3] ),
    .ZN(_07095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12380_ (.A1(_06969_),
    .A2(_07088_),
    .B(_07095_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12381_ (.A1(_07094_),
    .A2(\register_file[24][4] ),
    .ZN(_07096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12382_ (.A1(_06972_),
    .A2(_07088_),
    .B(_07096_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12383_ (.I(_07089_),
    .Z(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12384_ (.I(_07097_),
    .Z(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12385_ (.A1(_07094_),
    .A2(\register_file[24][5] ),
    .ZN(_07099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12386_ (.A1(_06974_),
    .A2(_07098_),
    .B(_07099_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12387_ (.A1(_07094_),
    .A2(\register_file[24][6] ),
    .ZN(_07100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12388_ (.A1(_06978_),
    .A2(_07098_),
    .B(_07100_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12389_ (.A1(_07094_),
    .A2(\register_file[24][7] ),
    .ZN(_07101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12390_ (.A1(_06980_),
    .A2(_07098_),
    .B(_07101_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12391_ (.I(_07089_),
    .Z(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12392_ (.A1(_07102_),
    .A2(\register_file[24][8] ),
    .ZN(_07103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12393_ (.A1(_06982_),
    .A2(_07098_),
    .B(_07103_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12394_ (.A1(_07102_),
    .A2(\register_file[24][9] ),
    .ZN(_07104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12395_ (.A1(_06985_),
    .A2(_07098_),
    .B(_07104_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12396_ (.I(_07097_),
    .Z(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12397_ (.A1(_07102_),
    .A2(\register_file[24][10] ),
    .ZN(_07106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12398_ (.A1(_06987_),
    .A2(_07105_),
    .B(_07106_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12399_ (.A1(_07102_),
    .A2(\register_file[24][11] ),
    .ZN(_07107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12400_ (.A1(_06990_),
    .A2(_07105_),
    .B(_07107_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12401_ (.A1(_07102_),
    .A2(\register_file[24][12] ),
    .ZN(_07108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12402_ (.A1(_06992_),
    .A2(_07105_),
    .B(_07108_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12403_ (.I(_07089_),
    .Z(_07109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12404_ (.A1(_07109_),
    .A2(\register_file[24][13] ),
    .ZN(_07110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12405_ (.A1(_06994_),
    .A2(_07105_),
    .B(_07110_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12406_ (.A1(_07109_),
    .A2(\register_file[24][14] ),
    .ZN(_07111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12407_ (.A1(_06997_),
    .A2(_07105_),
    .B(_07111_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12408_ (.I(_07097_),
    .Z(_07112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12409_ (.A1(_07109_),
    .A2(\register_file[24][15] ),
    .ZN(_07113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12410_ (.A1(_06999_),
    .A2(_07112_),
    .B(_07113_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12411_ (.A1(_07109_),
    .A2(\register_file[24][16] ),
    .ZN(_07114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12412_ (.A1(_07002_),
    .A2(_07112_),
    .B(_07114_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12413_ (.A1(_07109_),
    .A2(\register_file[24][17] ),
    .ZN(_07115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12414_ (.A1(_07004_),
    .A2(_07112_),
    .B(_07115_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12415_ (.I(_07086_),
    .Z(_07116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12416_ (.A1(_07116_),
    .A2(\register_file[24][18] ),
    .ZN(_07117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12417_ (.A1(_07006_),
    .A2(_07112_),
    .B(_07117_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12418_ (.A1(_07116_),
    .A2(\register_file[24][19] ),
    .ZN(_07118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12419_ (.A1(_07009_),
    .A2(_07112_),
    .B(_07118_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12420_ (.I(_07097_),
    .Z(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12421_ (.A1(_07116_),
    .A2(\register_file[24][20] ),
    .ZN(_07120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12422_ (.A1(_07011_),
    .A2(_07119_),
    .B(_07120_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12423_ (.A1(_07116_),
    .A2(\register_file[24][21] ),
    .ZN(_07121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12424_ (.A1(_07014_),
    .A2(_07119_),
    .B(_07121_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12425_ (.A1(_07116_),
    .A2(\register_file[24][22] ),
    .ZN(_07122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12426_ (.A1(_07016_),
    .A2(_07119_),
    .B(_07122_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12427_ (.I(_07086_),
    .Z(_07123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12428_ (.A1(_07123_),
    .A2(\register_file[24][23] ),
    .ZN(_07124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12429_ (.A1(_07018_),
    .A2(_07119_),
    .B(_07124_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12430_ (.A1(_07123_),
    .A2(\register_file[24][24] ),
    .ZN(_07125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12431_ (.A1(_07021_),
    .A2(_07119_),
    .B(_07125_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12432_ (.I(_07097_),
    .Z(_07126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12433_ (.A1(_07123_),
    .A2(\register_file[24][25] ),
    .ZN(_07127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12434_ (.A1(_07023_),
    .A2(_07126_),
    .B(_07127_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12435_ (.A1(_07123_),
    .A2(\register_file[24][26] ),
    .ZN(_07128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12436_ (.A1(_07026_),
    .A2(_07126_),
    .B(_07128_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12437_ (.A1(_07123_),
    .A2(\register_file[24][27] ),
    .ZN(_07129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12438_ (.A1(_07028_),
    .A2(_07126_),
    .B(_07129_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12439_ (.A1(_07087_),
    .A2(\register_file[24][28] ),
    .ZN(_07130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12440_ (.A1(_07030_),
    .A2(_07126_),
    .B(_07130_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12441_ (.A1(_07087_),
    .A2(\register_file[24][29] ),
    .ZN(_07131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12442_ (.A1(_07032_),
    .A2(_07126_),
    .B(_07131_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12443_ (.A1(_07087_),
    .A2(\register_file[24][30] ),
    .ZN(_07132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12444_ (.A1(_07034_),
    .A2(_07090_),
    .B(_07132_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12445_ (.A1(_07087_),
    .A2(\register_file[24][31] ),
    .ZN(_07133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12446_ (.A1(_07036_),
    .A2(_07090_),
    .B(_07133_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12447_ (.A1(_06265_),
    .A2(_03991_),
    .ZN(_07134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12448_ (.I(_07134_),
    .Z(_07135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12449_ (.I(_07135_),
    .Z(_07136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12450_ (.I(_07134_),
    .Z(_07137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12451_ (.I(_07137_),
    .Z(_07138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12452_ (.A1(_07138_),
    .A2(\register_file[23][0] ),
    .ZN(_07139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12453_ (.A1(_06958_),
    .A2(_07136_),
    .B(_07139_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12454_ (.A1(_07138_),
    .A2(\register_file[23][1] ),
    .ZN(_07140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12455_ (.A1(_06965_),
    .A2(_07136_),
    .B(_07140_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12456_ (.A1(_07138_),
    .A2(\register_file[23][2] ),
    .ZN(_07141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12457_ (.A1(_06967_),
    .A2(_07136_),
    .B(_07141_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12458_ (.I(_07137_),
    .Z(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12459_ (.A1(_07142_),
    .A2(\register_file[23][3] ),
    .ZN(_07143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12460_ (.A1(_06969_),
    .A2(_07136_),
    .B(_07143_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12461_ (.A1(_07142_),
    .A2(\register_file[23][4] ),
    .ZN(_07144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12462_ (.A1(_06972_),
    .A2(_07136_),
    .B(_07144_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12463_ (.I(_07137_),
    .Z(_07145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12464_ (.I(_07145_),
    .Z(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12465_ (.A1(_07142_),
    .A2(\register_file[23][5] ),
    .ZN(_07147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12466_ (.A1(_06974_),
    .A2(_07146_),
    .B(_07147_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12467_ (.A1(_07142_),
    .A2(\register_file[23][6] ),
    .ZN(_07148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12468_ (.A1(_06978_),
    .A2(_07146_),
    .B(_07148_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12469_ (.A1(_07142_),
    .A2(\register_file[23][7] ),
    .ZN(_07149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12470_ (.A1(_06980_),
    .A2(_07146_),
    .B(_07149_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12471_ (.I(_07137_),
    .Z(_07150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12472_ (.A1(_07150_),
    .A2(\register_file[23][8] ),
    .ZN(_07151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12473_ (.A1(_06982_),
    .A2(_07146_),
    .B(_07151_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12474_ (.A1(_07150_),
    .A2(\register_file[23][9] ),
    .ZN(_07152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12475_ (.A1(_06985_),
    .A2(_07146_),
    .B(_07152_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12476_ (.I(_07145_),
    .Z(_07153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12477_ (.A1(_07150_),
    .A2(\register_file[23][10] ),
    .ZN(_07154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12478_ (.A1(_06987_),
    .A2(_07153_),
    .B(_07154_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12479_ (.A1(_07150_),
    .A2(\register_file[23][11] ),
    .ZN(_07155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12480_ (.A1(_06990_),
    .A2(_07153_),
    .B(_07155_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12481_ (.A1(_07150_),
    .A2(\register_file[23][12] ),
    .ZN(_07156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12482_ (.A1(_06992_),
    .A2(_07153_),
    .B(_07156_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12483_ (.I(_07137_),
    .Z(_07157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12484_ (.A1(_07157_),
    .A2(\register_file[23][13] ),
    .ZN(_07158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12485_ (.A1(_06994_),
    .A2(_07153_),
    .B(_07158_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12486_ (.A1(_07157_),
    .A2(\register_file[23][14] ),
    .ZN(_07159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12487_ (.A1(_06997_),
    .A2(_07153_),
    .B(_07159_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12488_ (.I(_07145_),
    .Z(_07160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12489_ (.A1(_07157_),
    .A2(\register_file[23][15] ),
    .ZN(_07161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12490_ (.A1(_06999_),
    .A2(_07160_),
    .B(_07161_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12491_ (.A1(_07157_),
    .A2(\register_file[23][16] ),
    .ZN(_07162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12492_ (.A1(_07002_),
    .A2(_07160_),
    .B(_07162_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12493_ (.A1(_07157_),
    .A2(\register_file[23][17] ),
    .ZN(_07163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12494_ (.A1(_07004_),
    .A2(_07160_),
    .B(_07163_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12495_ (.I(_07134_),
    .Z(_07164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12496_ (.A1(_07164_),
    .A2(\register_file[23][18] ),
    .ZN(_07165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12497_ (.A1(_07006_),
    .A2(_07160_),
    .B(_07165_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12498_ (.A1(_07164_),
    .A2(\register_file[23][19] ),
    .ZN(_07166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12499_ (.A1(_07009_),
    .A2(_07160_),
    .B(_07166_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12500_ (.I(_07145_),
    .Z(_07167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12501_ (.A1(_07164_),
    .A2(\register_file[23][20] ),
    .ZN(_07168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12502_ (.A1(_07011_),
    .A2(_07167_),
    .B(_07168_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12503_ (.A1(_07164_),
    .A2(\register_file[23][21] ),
    .ZN(_07169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12504_ (.A1(_07014_),
    .A2(_07167_),
    .B(_07169_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12505_ (.A1(_07164_),
    .A2(\register_file[23][22] ),
    .ZN(_07170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12506_ (.A1(_07016_),
    .A2(_07167_),
    .B(_07170_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12507_ (.I(_07134_),
    .Z(_07171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12508_ (.A1(_07171_),
    .A2(\register_file[23][23] ),
    .ZN(_07172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12509_ (.A1(_07018_),
    .A2(_07167_),
    .B(_07172_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12510_ (.A1(_07171_),
    .A2(\register_file[23][24] ),
    .ZN(_07173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12511_ (.A1(_07021_),
    .A2(_07167_),
    .B(_07173_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12512_ (.I(_07145_),
    .Z(_07174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12513_ (.A1(_07171_),
    .A2(\register_file[23][25] ),
    .ZN(_07175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12514_ (.A1(_07023_),
    .A2(_07174_),
    .B(_07175_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12515_ (.A1(_07171_),
    .A2(\register_file[23][26] ),
    .ZN(_07176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12516_ (.A1(_07026_),
    .A2(_07174_),
    .B(_07176_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12517_ (.A1(_07171_),
    .A2(\register_file[23][27] ),
    .ZN(_07177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12518_ (.A1(_07028_),
    .A2(_07174_),
    .B(_07177_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12519_ (.A1(_07135_),
    .A2(\register_file[23][28] ),
    .ZN(_07178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12520_ (.A1(_07030_),
    .A2(_07174_),
    .B(_07178_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12521_ (.A1(_07135_),
    .A2(\register_file[23][29] ),
    .ZN(_07179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12522_ (.A1(_07032_),
    .A2(_07174_),
    .B(_07179_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12523_ (.A1(_07135_),
    .A2(\register_file[23][30] ),
    .ZN(_07180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12524_ (.A1(_07034_),
    .A2(_07138_),
    .B(_07180_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12525_ (.A1(_07135_),
    .A2(\register_file[23][31] ),
    .ZN(_07181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12526_ (.A1(_07036_),
    .A2(_07138_),
    .B(_07181_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12527_ (.A1(_06023_),
    .A2(_03991_),
    .ZN(_07182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12528_ (.I(_07182_),
    .Z(_07183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12529_ (.I(_07183_),
    .Z(_07184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12530_ (.I(_07182_),
    .Z(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12531_ (.I(_07185_),
    .Z(_07186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12532_ (.A1(_07186_),
    .A2(\register_file[22][0] ),
    .ZN(_07187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12533_ (.A1(_06958_),
    .A2(_07184_),
    .B(_07187_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12534_ (.A1(_07186_),
    .A2(\register_file[22][1] ),
    .ZN(_07188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12535_ (.A1(_06965_),
    .A2(_07184_),
    .B(_07188_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12536_ (.A1(_07186_),
    .A2(\register_file[22][2] ),
    .ZN(_07189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12537_ (.A1(_06967_),
    .A2(_07184_),
    .B(_07189_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12538_ (.I(_07185_),
    .Z(_07190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12539_ (.A1(_07190_),
    .A2(\register_file[22][3] ),
    .ZN(_07191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12540_ (.A1(_06969_),
    .A2(_07184_),
    .B(_07191_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12541_ (.A1(_07190_),
    .A2(\register_file[22][4] ),
    .ZN(_07192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12542_ (.A1(_06972_),
    .A2(_07184_),
    .B(_07192_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12543_ (.I(_07185_),
    .Z(_07193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12544_ (.I(_07193_),
    .Z(_07194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12545_ (.A1(_07190_),
    .A2(\register_file[22][5] ),
    .ZN(_07195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12546_ (.A1(_06974_),
    .A2(_07194_),
    .B(_07195_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12547_ (.A1(_07190_),
    .A2(\register_file[22][6] ),
    .ZN(_07196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12548_ (.A1(_06978_),
    .A2(_07194_),
    .B(_07196_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12549_ (.A1(_07190_),
    .A2(\register_file[22][7] ),
    .ZN(_07197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12550_ (.A1(_06980_),
    .A2(_07194_),
    .B(_07197_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12551_ (.I(_07185_),
    .Z(_07198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12552_ (.A1(_07198_),
    .A2(\register_file[22][8] ),
    .ZN(_07199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12553_ (.A1(_06982_),
    .A2(_07194_),
    .B(_07199_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12554_ (.A1(_07198_),
    .A2(\register_file[22][9] ),
    .ZN(_07200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12555_ (.A1(_06985_),
    .A2(_07194_),
    .B(_07200_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12556_ (.I(_07193_),
    .Z(_07201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12557_ (.A1(_07198_),
    .A2(\register_file[22][10] ),
    .ZN(_07202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12558_ (.A1(_06987_),
    .A2(_07201_),
    .B(_07202_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12559_ (.A1(_07198_),
    .A2(\register_file[22][11] ),
    .ZN(_07203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12560_ (.A1(_06990_),
    .A2(_07201_),
    .B(_07203_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12561_ (.A1(_07198_),
    .A2(\register_file[22][12] ),
    .ZN(_07204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12562_ (.A1(_06992_),
    .A2(_07201_),
    .B(_07204_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12563_ (.I(_07185_),
    .Z(_07205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12564_ (.A1(_07205_),
    .A2(\register_file[22][13] ),
    .ZN(_07206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12565_ (.A1(_06994_),
    .A2(_07201_),
    .B(_07206_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12566_ (.A1(_07205_),
    .A2(\register_file[22][14] ),
    .ZN(_07207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12567_ (.A1(_06997_),
    .A2(_07201_),
    .B(_07207_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12568_ (.I(_07193_),
    .Z(_07208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12569_ (.A1(_07205_),
    .A2(\register_file[22][15] ),
    .ZN(_07209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12570_ (.A1(_06999_),
    .A2(_07208_),
    .B(_07209_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12571_ (.A1(_07205_),
    .A2(\register_file[22][16] ),
    .ZN(_07210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12572_ (.A1(_07002_),
    .A2(_07208_),
    .B(_07210_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12573_ (.A1(_07205_),
    .A2(\register_file[22][17] ),
    .ZN(_07211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12574_ (.A1(_07004_),
    .A2(_07208_),
    .B(_07211_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12575_ (.I(_07182_),
    .Z(_07212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12576_ (.A1(_07212_),
    .A2(\register_file[22][18] ),
    .ZN(_07213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12577_ (.A1(_07006_),
    .A2(_07208_),
    .B(_07213_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12578_ (.A1(_07212_),
    .A2(\register_file[22][19] ),
    .ZN(_07214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12579_ (.A1(_07009_),
    .A2(_07208_),
    .B(_07214_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12580_ (.I(_07193_),
    .Z(_07215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12581_ (.A1(_07212_),
    .A2(\register_file[22][20] ),
    .ZN(_07216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12582_ (.A1(_07011_),
    .A2(_07215_),
    .B(_07216_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12583_ (.A1(_07212_),
    .A2(\register_file[22][21] ),
    .ZN(_07217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12584_ (.A1(_07014_),
    .A2(_07215_),
    .B(_07217_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12585_ (.A1(_07212_),
    .A2(\register_file[22][22] ),
    .ZN(_07218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12586_ (.A1(_07016_),
    .A2(_07215_),
    .B(_07218_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12587_ (.I(_07182_),
    .Z(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12588_ (.A1(_07219_),
    .A2(\register_file[22][23] ),
    .ZN(_07220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12589_ (.A1(_07018_),
    .A2(_07215_),
    .B(_07220_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12590_ (.A1(_07219_),
    .A2(\register_file[22][24] ),
    .ZN(_07221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12591_ (.A1(_07021_),
    .A2(_07215_),
    .B(_07221_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12592_ (.I(_07193_),
    .Z(_07222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12593_ (.A1(_07219_),
    .A2(\register_file[22][25] ),
    .ZN(_07223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12594_ (.A1(_07023_),
    .A2(_07222_),
    .B(_07223_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12595_ (.A1(_07219_),
    .A2(\register_file[22][26] ),
    .ZN(_07224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12596_ (.A1(_07026_),
    .A2(_07222_),
    .B(_07224_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12597_ (.A1(_07219_),
    .A2(\register_file[22][27] ),
    .ZN(_07225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12598_ (.A1(_07028_),
    .A2(_07222_),
    .B(_07225_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12599_ (.A1(_07183_),
    .A2(\register_file[22][28] ),
    .ZN(_07226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12600_ (.A1(_07030_),
    .A2(_07222_),
    .B(_07226_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12601_ (.A1(_07183_),
    .A2(\register_file[22][29] ),
    .ZN(_07227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12602_ (.A1(_07032_),
    .A2(_07222_),
    .B(_07227_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12603_ (.A1(_07183_),
    .A2(\register_file[22][30] ),
    .ZN(_07228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12604_ (.A1(_07034_),
    .A2(_07186_),
    .B(_07228_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12605_ (.A1(_07183_),
    .A2(\register_file[22][31] ),
    .ZN(_07229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12606_ (.A1(_07036_),
    .A2(_07186_),
    .B(_07229_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12607_ (.I(_06020_),
    .Z(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12608_ (.A1(_06317_),
    .A2(_03836_),
    .ZN(_07231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12609_ (.I(_07231_),
    .Z(_07232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12610_ (.I(_07232_),
    .Z(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12611_ (.I(_07231_),
    .Z(_07234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12612_ (.I(_07234_),
    .Z(_07235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12613_ (.A1(_07235_),
    .A2(\register_file[21][0] ),
    .ZN(_07236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12614_ (.A1(_07230_),
    .A2(_07233_),
    .B(_07236_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12615_ (.I(_06032_),
    .Z(_07237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12616_ (.A1(_07235_),
    .A2(\register_file[21][1] ),
    .ZN(_07238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12617_ (.A1(_07237_),
    .A2(_07233_),
    .B(_07238_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12618_ (.I(_06036_),
    .Z(_07239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12619_ (.A1(_07235_),
    .A2(\register_file[21][2] ),
    .ZN(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12620_ (.A1(_07239_),
    .A2(_07233_),
    .B(_07240_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12621_ (.I(_06040_),
    .Z(_07241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12622_ (.I(_07234_),
    .Z(_07242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12623_ (.A1(_07242_),
    .A2(\register_file[21][3] ),
    .ZN(_07243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12624_ (.A1(_07241_),
    .A2(_07233_),
    .B(_07243_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12625_ (.I(_06045_),
    .Z(_07244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12626_ (.A1(_07242_),
    .A2(\register_file[21][4] ),
    .ZN(_07245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12627_ (.A1(_07244_),
    .A2(_07233_),
    .B(_07245_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12628_ (.I(_06049_),
    .Z(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _12629_ (.I(_07234_),
    .Z(_07247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12630_ (.I(_07247_),
    .Z(_07248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12631_ (.A1(_07242_),
    .A2(\register_file[21][5] ),
    .ZN(_07249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12632_ (.A1(_07246_),
    .A2(_07248_),
    .B(_07249_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12633_ (.I(_06055_),
    .Z(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12634_ (.A1(_07242_),
    .A2(\register_file[21][6] ),
    .ZN(_07251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12635_ (.A1(_07250_),
    .A2(_07248_),
    .B(_07251_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12636_ (.I(_06059_),
    .Z(_07252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12637_ (.A1(_07242_),
    .A2(\register_file[21][7] ),
    .ZN(_07253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12638_ (.A1(_07252_),
    .A2(_07248_),
    .B(_07253_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12639_ (.I(_06063_),
    .Z(_07254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12640_ (.I(_07234_),
    .Z(_07255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12641_ (.A1(_07255_),
    .A2(\register_file[21][8] ),
    .ZN(_07256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12642_ (.A1(_07254_),
    .A2(_07248_),
    .B(_07256_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12643_ (.I(_06068_),
    .Z(_07257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12644_ (.A1(_07255_),
    .A2(\register_file[21][9] ),
    .ZN(_07258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12645_ (.A1(_07257_),
    .A2(_07248_),
    .B(_07258_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12646_ (.I(_06072_),
    .Z(_07259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12647_ (.I(_07247_),
    .Z(_07260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12648_ (.A1(_07255_),
    .A2(\register_file[21][10] ),
    .ZN(_07261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12649_ (.A1(_07259_),
    .A2(_07260_),
    .B(_07261_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12650_ (.I(_06077_),
    .Z(_07262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12651_ (.A1(_07255_),
    .A2(\register_file[21][11] ),
    .ZN(_07263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12652_ (.A1(_07262_),
    .A2(_07260_),
    .B(_07263_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12653_ (.I(_06081_),
    .Z(_07264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12654_ (.A1(_07255_),
    .A2(\register_file[21][12] ),
    .ZN(_07265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12655_ (.A1(_07264_),
    .A2(_07260_),
    .B(_07265_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12656_ (.I(_06085_),
    .Z(_07266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12657_ (.I(_07234_),
    .Z(_07267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12658_ (.A1(_07267_),
    .A2(\register_file[21][13] ),
    .ZN(_07268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12659_ (.A1(_07266_),
    .A2(_07260_),
    .B(_07268_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12660_ (.I(_06090_),
    .Z(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12661_ (.A1(_07267_),
    .A2(\register_file[21][14] ),
    .ZN(_07270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12662_ (.A1(_07269_),
    .A2(_07260_),
    .B(_07270_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12663_ (.I(_06094_),
    .Z(_07271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12664_ (.I(_07247_),
    .Z(_07272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12665_ (.A1(_07267_),
    .A2(\register_file[21][15] ),
    .ZN(_07273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12666_ (.A1(_07271_),
    .A2(_07272_),
    .B(_07273_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12667_ (.I(_06099_),
    .Z(_07274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12668_ (.A1(_07267_),
    .A2(\register_file[21][16] ),
    .ZN(_07275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12669_ (.A1(_07274_),
    .A2(_07272_),
    .B(_07275_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12670_ (.I(_06103_),
    .Z(_07276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12671_ (.A1(_07267_),
    .A2(\register_file[21][17] ),
    .ZN(_07277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12672_ (.A1(_07276_),
    .A2(_07272_),
    .B(_07277_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12673_ (.I(_06107_),
    .Z(_07278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12674_ (.I(_07231_),
    .Z(_07279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12675_ (.A1(_07279_),
    .A2(\register_file[21][18] ),
    .ZN(_07280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12676_ (.A1(_07278_),
    .A2(_07272_),
    .B(_07280_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12677_ (.I(_06112_),
    .Z(_07281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12678_ (.A1(_07279_),
    .A2(\register_file[21][19] ),
    .ZN(_07282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12679_ (.A1(_07281_),
    .A2(_07272_),
    .B(_07282_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12680_ (.I(_06116_),
    .Z(_07283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12681_ (.I(_07247_),
    .Z(_07284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12682_ (.A1(_07279_),
    .A2(\register_file[21][20] ),
    .ZN(_07285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12683_ (.A1(_07283_),
    .A2(_07284_),
    .B(_07285_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12684_ (.I(_06121_),
    .Z(_07286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12685_ (.A1(_07279_),
    .A2(\register_file[21][21] ),
    .ZN(_07287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12686_ (.A1(_07286_),
    .A2(_07284_),
    .B(_07287_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12687_ (.I(_06125_),
    .Z(_07288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12688_ (.A1(_07279_),
    .A2(\register_file[21][22] ),
    .ZN(_07289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12689_ (.A1(_07288_),
    .A2(_07284_),
    .B(_07289_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12690_ (.I(_06129_),
    .Z(_07290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12691_ (.I(_07231_),
    .Z(_07291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12692_ (.A1(_07291_),
    .A2(\register_file[21][23] ),
    .ZN(_07292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12693_ (.A1(_07290_),
    .A2(_07284_),
    .B(_07292_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12694_ (.I(_06134_),
    .Z(_07293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12695_ (.A1(_07291_),
    .A2(\register_file[21][24] ),
    .ZN(_07294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12696_ (.A1(_07293_),
    .A2(_07284_),
    .B(_07294_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12697_ (.I(_06138_),
    .Z(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12698_ (.I(_07247_),
    .Z(_07296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12699_ (.A1(_07291_),
    .A2(\register_file[21][25] ),
    .ZN(_07297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12700_ (.A1(_07295_),
    .A2(_07296_),
    .B(_07297_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12701_ (.I(_06143_),
    .Z(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12702_ (.A1(_07291_),
    .A2(\register_file[21][26] ),
    .ZN(_07299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12703_ (.A1(_07298_),
    .A2(_07296_),
    .B(_07299_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12704_ (.I(_06147_),
    .Z(_07300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12705_ (.A1(_07291_),
    .A2(\register_file[21][27] ),
    .ZN(_07301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12706_ (.A1(_07300_),
    .A2(_07296_),
    .B(_07301_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12707_ (.I(_06151_),
    .Z(_07302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12708_ (.A1(_07232_),
    .A2(\register_file[21][28] ),
    .ZN(_07303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12709_ (.A1(_07302_),
    .A2(_07296_),
    .B(_07303_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12710_ (.I(_06155_),
    .Z(_07304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12711_ (.A1(_07232_),
    .A2(\register_file[21][29] ),
    .ZN(_07305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12712_ (.A1(_07304_),
    .A2(_07296_),
    .B(_07305_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12713_ (.I(_06159_),
    .Z(_07306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12714_ (.A1(_07232_),
    .A2(\register_file[21][30] ),
    .ZN(_07307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12715_ (.A1(_07306_),
    .A2(_07235_),
    .B(_07307_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12716_ (.I(_06163_),
    .Z(_07308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12717_ (.A1(_07232_),
    .A2(\register_file[21][31] ),
    .ZN(_07309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12718_ (.A1(_07308_),
    .A2(_07235_),
    .B(_07309_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12719_ (.A1(_06216_),
    .A2(_03836_),
    .ZN(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12720_ (.I(_07310_),
    .Z(_07311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12721_ (.I(_07311_),
    .Z(_07312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12722_ (.I(_07310_),
    .Z(_07313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12723_ (.I(_07313_),
    .Z(_07314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12724_ (.A1(_07314_),
    .A2(\register_file[20][0] ),
    .ZN(_07315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12725_ (.A1(_07230_),
    .A2(_07312_),
    .B(_07315_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12726_ (.A1(_07314_),
    .A2(\register_file[20][1] ),
    .ZN(_07316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12727_ (.A1(_07237_),
    .A2(_07312_),
    .B(_07316_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12728_ (.A1(_07314_),
    .A2(\register_file[20][2] ),
    .ZN(_07317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12729_ (.A1(_07239_),
    .A2(_07312_),
    .B(_07317_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12730_ (.I(_07313_),
    .Z(_07318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12731_ (.A1(_07318_),
    .A2(\register_file[20][3] ),
    .ZN(_07319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12732_ (.A1(_07241_),
    .A2(_07312_),
    .B(_07319_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12733_ (.A1(_07318_),
    .A2(\register_file[20][4] ),
    .ZN(_07320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12734_ (.A1(_07244_),
    .A2(_07312_),
    .B(_07320_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12735_ (.I(_07313_),
    .Z(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12736_ (.I(_07321_),
    .Z(_07322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12737_ (.A1(_07318_),
    .A2(\register_file[20][5] ),
    .ZN(_07323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12738_ (.A1(_07246_),
    .A2(_07322_),
    .B(_07323_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12739_ (.A1(_07318_),
    .A2(\register_file[20][6] ),
    .ZN(_07324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12740_ (.A1(_07250_),
    .A2(_07322_),
    .B(_07324_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12741_ (.A1(_07318_),
    .A2(\register_file[20][7] ),
    .ZN(_07325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12742_ (.A1(_07252_),
    .A2(_07322_),
    .B(_07325_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12743_ (.I(_07313_),
    .Z(_07326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12744_ (.A1(_07326_),
    .A2(\register_file[20][8] ),
    .ZN(_07327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12745_ (.A1(_07254_),
    .A2(_07322_),
    .B(_07327_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12746_ (.A1(_07326_),
    .A2(\register_file[20][9] ),
    .ZN(_07328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12747_ (.A1(_07257_),
    .A2(_07322_),
    .B(_07328_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12748_ (.I(_07321_),
    .Z(_07329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12749_ (.A1(_07326_),
    .A2(\register_file[20][10] ),
    .ZN(_07330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12750_ (.A1(_07259_),
    .A2(_07329_),
    .B(_07330_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12751_ (.A1(_07326_),
    .A2(\register_file[20][11] ),
    .ZN(_07331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12752_ (.A1(_07262_),
    .A2(_07329_),
    .B(_07331_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12753_ (.A1(_07326_),
    .A2(\register_file[20][12] ),
    .ZN(_07332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12754_ (.A1(_07264_),
    .A2(_07329_),
    .B(_07332_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12755_ (.I(_07313_),
    .Z(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12756_ (.A1(_07333_),
    .A2(\register_file[20][13] ),
    .ZN(_07334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12757_ (.A1(_07266_),
    .A2(_07329_),
    .B(_07334_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12758_ (.A1(_07333_),
    .A2(\register_file[20][14] ),
    .ZN(_07335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12759_ (.A1(_07269_),
    .A2(_07329_),
    .B(_07335_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12760_ (.I(_07321_),
    .Z(_07336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12761_ (.A1(_07333_),
    .A2(\register_file[20][15] ),
    .ZN(_07337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12762_ (.A1(_07271_),
    .A2(_07336_),
    .B(_07337_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12763_ (.A1(_07333_),
    .A2(\register_file[20][16] ),
    .ZN(_07338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12764_ (.A1(_07274_),
    .A2(_07336_),
    .B(_07338_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12765_ (.A1(_07333_),
    .A2(\register_file[20][17] ),
    .ZN(_07339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12766_ (.A1(_07276_),
    .A2(_07336_),
    .B(_07339_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12767_ (.I(_07310_),
    .Z(_07340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12768_ (.A1(_07340_),
    .A2(\register_file[20][18] ),
    .ZN(_07341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12769_ (.A1(_07278_),
    .A2(_07336_),
    .B(_07341_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12770_ (.A1(_07340_),
    .A2(\register_file[20][19] ),
    .ZN(_07342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12771_ (.A1(_07281_),
    .A2(_07336_),
    .B(_07342_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12772_ (.I(_07321_),
    .Z(_07343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12773_ (.A1(_07340_),
    .A2(\register_file[20][20] ),
    .ZN(_07344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12774_ (.A1(_07283_),
    .A2(_07343_),
    .B(_07344_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12775_ (.A1(_07340_),
    .A2(\register_file[20][21] ),
    .ZN(_07345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12776_ (.A1(_07286_),
    .A2(_07343_),
    .B(_07345_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12777_ (.A1(_07340_),
    .A2(\register_file[20][22] ),
    .ZN(_07346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12778_ (.A1(_07288_),
    .A2(_07343_),
    .B(_07346_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12779_ (.I(_07310_),
    .Z(_07347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12780_ (.A1(_07347_),
    .A2(\register_file[20][23] ),
    .ZN(_07348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12781_ (.A1(_07290_),
    .A2(_07343_),
    .B(_07348_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12782_ (.A1(_07347_),
    .A2(\register_file[20][24] ),
    .ZN(_07349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12783_ (.A1(_07293_),
    .A2(_07343_),
    .B(_07349_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12784_ (.I(_07321_),
    .Z(_07350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12785_ (.A1(_07347_),
    .A2(\register_file[20][25] ),
    .ZN(_07351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12786_ (.A1(_07295_),
    .A2(_07350_),
    .B(_07351_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12787_ (.A1(_07347_),
    .A2(\register_file[20][26] ),
    .ZN(_07352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12788_ (.A1(_07298_),
    .A2(_07350_),
    .B(_07352_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12789_ (.A1(_07347_),
    .A2(\register_file[20][27] ),
    .ZN(_07353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12790_ (.A1(_07300_),
    .A2(_07350_),
    .B(_07353_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12791_ (.A1(_07311_),
    .A2(\register_file[20][28] ),
    .ZN(_07354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12792_ (.A1(_07302_),
    .A2(_07350_),
    .B(_07354_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12793_ (.A1(_07311_),
    .A2(\register_file[20][29] ),
    .ZN(_07355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12794_ (.A1(_07304_),
    .A2(_07350_),
    .B(_07355_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12795_ (.A1(_07311_),
    .A2(\register_file[20][30] ),
    .ZN(_07356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12796_ (.A1(_07306_),
    .A2(_07314_),
    .B(_07356_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12797_ (.A1(_07311_),
    .A2(\register_file[20][31] ),
    .ZN(_07357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12798_ (.A1(_07308_),
    .A2(_07314_),
    .B(_07357_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12799_ (.A1(_06317_),
    .A2(_03927_),
    .ZN(_07358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12800_ (.I(_07358_),
    .Z(_07359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12801_ (.I(_07359_),
    .Z(_07360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12802_ (.I(_07358_),
    .Z(_07361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12803_ (.I(_07361_),
    .Z(_07362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12804_ (.A1(_07362_),
    .A2(\register_file[1][0] ),
    .ZN(_07363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12805_ (.A1(_07230_),
    .A2(_07360_),
    .B(_07363_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12806_ (.A1(_07362_),
    .A2(\register_file[1][1] ),
    .ZN(_07364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12807_ (.A1(_07237_),
    .A2(_07360_),
    .B(_07364_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12808_ (.A1(_07362_),
    .A2(\register_file[1][2] ),
    .ZN(_07365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12809_ (.A1(_07239_),
    .A2(_07360_),
    .B(_07365_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12810_ (.I(_07361_),
    .Z(_07366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12811_ (.A1(_07366_),
    .A2(\register_file[1][3] ),
    .ZN(_07367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12812_ (.A1(_07241_),
    .A2(_07360_),
    .B(_07367_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12813_ (.A1(_07366_),
    .A2(\register_file[1][4] ),
    .ZN(_07368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12814_ (.A1(_07244_),
    .A2(_07360_),
    .B(_07368_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12815_ (.I(_07361_),
    .Z(_07369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12816_ (.I(_07369_),
    .Z(_07370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12817_ (.A1(_07366_),
    .A2(\register_file[1][5] ),
    .ZN(_07371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12818_ (.A1(_07246_),
    .A2(_07370_),
    .B(_07371_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12819_ (.A1(_07366_),
    .A2(\register_file[1][6] ),
    .ZN(_07372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12820_ (.A1(_07250_),
    .A2(_07370_),
    .B(_07372_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12821_ (.A1(_07366_),
    .A2(\register_file[1][7] ),
    .ZN(_07373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12822_ (.A1(_07252_),
    .A2(_07370_),
    .B(_07373_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12823_ (.I(_07361_),
    .Z(_07374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12824_ (.A1(_07374_),
    .A2(\register_file[1][8] ),
    .ZN(_07375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12825_ (.A1(_07254_),
    .A2(_07370_),
    .B(_07375_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12826_ (.A1(_07374_),
    .A2(\register_file[1][9] ),
    .ZN(_07376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12827_ (.A1(_07257_),
    .A2(_07370_),
    .B(_07376_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12828_ (.I(_07369_),
    .Z(_07377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12829_ (.A1(_07374_),
    .A2(\register_file[1][10] ),
    .ZN(_07378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12830_ (.A1(_07259_),
    .A2(_07377_),
    .B(_07378_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12831_ (.A1(_07374_),
    .A2(\register_file[1][11] ),
    .ZN(_07379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12832_ (.A1(_07262_),
    .A2(_07377_),
    .B(_07379_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12833_ (.A1(_07374_),
    .A2(\register_file[1][12] ),
    .ZN(_07380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12834_ (.A1(_07264_),
    .A2(_07377_),
    .B(_07380_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12835_ (.I(_07361_),
    .Z(_07381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12836_ (.A1(_07381_),
    .A2(\register_file[1][13] ),
    .ZN(_07382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12837_ (.A1(_07266_),
    .A2(_07377_),
    .B(_07382_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12838_ (.A1(_07381_),
    .A2(\register_file[1][14] ),
    .ZN(_07383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12839_ (.A1(_07269_),
    .A2(_07377_),
    .B(_07383_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12840_ (.I(_07369_),
    .Z(_07384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12841_ (.A1(_07381_),
    .A2(\register_file[1][15] ),
    .ZN(_07385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12842_ (.A1(_07271_),
    .A2(_07384_),
    .B(_07385_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12843_ (.A1(_07381_),
    .A2(\register_file[1][16] ),
    .ZN(_07386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12844_ (.A1(_07274_),
    .A2(_07384_),
    .B(_07386_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12845_ (.A1(_07381_),
    .A2(\register_file[1][17] ),
    .ZN(_07387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12846_ (.A1(_07276_),
    .A2(_07384_),
    .B(_07387_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12847_ (.I(_07358_),
    .Z(_07388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12848_ (.A1(_07388_),
    .A2(\register_file[1][18] ),
    .ZN(_07389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12849_ (.A1(_07278_),
    .A2(_07384_),
    .B(_07389_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12850_ (.A1(_07388_),
    .A2(\register_file[1][19] ),
    .ZN(_07390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12851_ (.A1(_07281_),
    .A2(_07384_),
    .B(_07390_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12852_ (.I(_07369_),
    .Z(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12853_ (.A1(_07388_),
    .A2(\register_file[1][20] ),
    .ZN(_07392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12854_ (.A1(_07283_),
    .A2(_07391_),
    .B(_07392_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12855_ (.A1(_07388_),
    .A2(\register_file[1][21] ),
    .ZN(_07393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12856_ (.A1(_07286_),
    .A2(_07391_),
    .B(_07393_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12857_ (.A1(_07388_),
    .A2(\register_file[1][22] ),
    .ZN(_07394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12858_ (.A1(_07288_),
    .A2(_07391_),
    .B(_07394_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12859_ (.I(_07358_),
    .Z(_07395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12860_ (.A1(_07395_),
    .A2(\register_file[1][23] ),
    .ZN(_07396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12861_ (.A1(_07290_),
    .A2(_07391_),
    .B(_07396_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12862_ (.A1(_07395_),
    .A2(\register_file[1][24] ),
    .ZN(_07397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12863_ (.A1(_07293_),
    .A2(_07391_),
    .B(_07397_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12864_ (.I(_07369_),
    .Z(_07398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12865_ (.A1(_07395_),
    .A2(\register_file[1][25] ),
    .ZN(_07399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12866_ (.A1(_07295_),
    .A2(_07398_),
    .B(_07399_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12867_ (.A1(_07395_),
    .A2(\register_file[1][26] ),
    .ZN(_07400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12868_ (.A1(_07298_),
    .A2(_07398_),
    .B(_07400_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12869_ (.A1(_07395_),
    .A2(\register_file[1][27] ),
    .ZN(_07401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12870_ (.A1(_07300_),
    .A2(_07398_),
    .B(_07401_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12871_ (.A1(_07359_),
    .A2(\register_file[1][28] ),
    .ZN(_07402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12872_ (.A1(_07302_),
    .A2(_07398_),
    .B(_07402_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12873_ (.A1(_07359_),
    .A2(\register_file[1][29] ),
    .ZN(_07403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12874_ (.A1(_07304_),
    .A2(_07398_),
    .B(_07403_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12875_ (.A1(_07359_),
    .A2(\register_file[1][30] ),
    .ZN(_07404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12876_ (.A1(_07306_),
    .A2(_07362_),
    .B(_07404_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12877_ (.A1(_07359_),
    .A2(\register_file[1][31] ),
    .ZN(_07405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12878_ (.A1(_07308_),
    .A2(_07362_),
    .B(_07405_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12879_ (.A1(_06023_),
    .A2(_03855_),
    .ZN(_07406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12880_ (.I(_07406_),
    .Z(_07407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12881_ (.I(_07407_),
    .Z(_07408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12882_ (.I(_07406_),
    .Z(_07409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12883_ (.I(_07409_),
    .Z(_07410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12884_ (.A1(_07410_),
    .A2(\register_file[18][0] ),
    .ZN(_07411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12885_ (.A1(_07230_),
    .A2(_07408_),
    .B(_07411_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12886_ (.A1(_07410_),
    .A2(\register_file[18][1] ),
    .ZN(_07412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12887_ (.A1(_07237_),
    .A2(_07408_),
    .B(_07412_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12888_ (.A1(_07410_),
    .A2(\register_file[18][2] ),
    .ZN(_07413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12889_ (.A1(_07239_),
    .A2(_07408_),
    .B(_07413_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12890_ (.I(_07409_),
    .Z(_07414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12891_ (.A1(_07414_),
    .A2(\register_file[18][3] ),
    .ZN(_07415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12892_ (.A1(_07241_),
    .A2(_07408_),
    .B(_07415_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12893_ (.A1(_07414_),
    .A2(\register_file[18][4] ),
    .ZN(_07416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12894_ (.A1(_07244_),
    .A2(_07408_),
    .B(_07416_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12895_ (.I(_07409_),
    .Z(_07417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12896_ (.I(_07417_),
    .Z(_07418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12897_ (.A1(_07414_),
    .A2(\register_file[18][5] ),
    .ZN(_07419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12898_ (.A1(_07246_),
    .A2(_07418_),
    .B(_07419_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12899_ (.A1(_07414_),
    .A2(\register_file[18][6] ),
    .ZN(_07420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12900_ (.A1(_07250_),
    .A2(_07418_),
    .B(_07420_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12901_ (.A1(_07414_),
    .A2(\register_file[18][7] ),
    .ZN(_07421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12902_ (.A1(_07252_),
    .A2(_07418_),
    .B(_07421_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12903_ (.I(_07409_),
    .Z(_07422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12904_ (.A1(_07422_),
    .A2(\register_file[18][8] ),
    .ZN(_07423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12905_ (.A1(_07254_),
    .A2(_07418_),
    .B(_07423_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12906_ (.A1(_07422_),
    .A2(\register_file[18][9] ),
    .ZN(_07424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12907_ (.A1(_07257_),
    .A2(_07418_),
    .B(_07424_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12908_ (.I(_07417_),
    .Z(_07425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12909_ (.A1(_07422_),
    .A2(\register_file[18][10] ),
    .ZN(_07426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12910_ (.A1(_07259_),
    .A2(_07425_),
    .B(_07426_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12911_ (.A1(_07422_),
    .A2(\register_file[18][11] ),
    .ZN(_07427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12912_ (.A1(_07262_),
    .A2(_07425_),
    .B(_07427_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12913_ (.A1(_07422_),
    .A2(\register_file[18][12] ),
    .ZN(_07428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12914_ (.A1(_07264_),
    .A2(_07425_),
    .B(_07428_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12915_ (.I(_07409_),
    .Z(_07429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12916_ (.A1(_07429_),
    .A2(\register_file[18][13] ),
    .ZN(_07430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12917_ (.A1(_07266_),
    .A2(_07425_),
    .B(_07430_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12918_ (.A1(_07429_),
    .A2(\register_file[18][14] ),
    .ZN(_07431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12919_ (.A1(_07269_),
    .A2(_07425_),
    .B(_07431_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12920_ (.I(_07417_),
    .Z(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12921_ (.A1(_07429_),
    .A2(\register_file[18][15] ),
    .ZN(_07433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12922_ (.A1(_07271_),
    .A2(_07432_),
    .B(_07433_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12923_ (.A1(_07429_),
    .A2(\register_file[18][16] ),
    .ZN(_07434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12924_ (.A1(_07274_),
    .A2(_07432_),
    .B(_07434_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12925_ (.A1(_07429_),
    .A2(\register_file[18][17] ),
    .ZN(_07435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12926_ (.A1(_07276_),
    .A2(_07432_),
    .B(_07435_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12927_ (.I(_07406_),
    .Z(_07436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12928_ (.A1(_07436_),
    .A2(\register_file[18][18] ),
    .ZN(_07437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12929_ (.A1(_07278_),
    .A2(_07432_),
    .B(_07437_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12930_ (.A1(_07436_),
    .A2(\register_file[18][19] ),
    .ZN(_07438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12931_ (.A1(_07281_),
    .A2(_07432_),
    .B(_07438_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12932_ (.I(_07417_),
    .Z(_07439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12933_ (.A1(_07436_),
    .A2(\register_file[18][20] ),
    .ZN(_07440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12934_ (.A1(_07283_),
    .A2(_07439_),
    .B(_07440_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12935_ (.A1(_07436_),
    .A2(\register_file[18][21] ),
    .ZN(_07441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12936_ (.A1(_07286_),
    .A2(_07439_),
    .B(_07441_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12937_ (.A1(_07436_),
    .A2(\register_file[18][22] ),
    .ZN(_07442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12938_ (.A1(_07288_),
    .A2(_07439_),
    .B(_07442_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12939_ (.I(_07406_),
    .Z(_07443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12940_ (.A1(_07443_),
    .A2(\register_file[18][23] ),
    .ZN(_07444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12941_ (.A1(_07290_),
    .A2(_07439_),
    .B(_07444_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12942_ (.A1(_07443_),
    .A2(\register_file[18][24] ),
    .ZN(_07445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12943_ (.A1(_07293_),
    .A2(_07439_),
    .B(_07445_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12944_ (.I(_07417_),
    .Z(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12945_ (.A1(_07443_),
    .A2(\register_file[18][25] ),
    .ZN(_07447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12946_ (.A1(_07295_),
    .A2(_07446_),
    .B(_07447_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12947_ (.A1(_07443_),
    .A2(\register_file[18][26] ),
    .ZN(_07448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12948_ (.A1(_07298_),
    .A2(_07446_),
    .B(_07448_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12949_ (.A1(_07443_),
    .A2(\register_file[18][27] ),
    .ZN(_07449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12950_ (.A1(_07300_),
    .A2(_07446_),
    .B(_07449_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12951_ (.A1(_07407_),
    .A2(\register_file[18][28] ),
    .ZN(_07450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12952_ (.A1(_07302_),
    .A2(_07446_),
    .B(_07450_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12953_ (.A1(_07407_),
    .A2(\register_file[18][29] ),
    .ZN(_07451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12954_ (.A1(_07304_),
    .A2(_07446_),
    .B(_07451_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12955_ (.A1(_07407_),
    .A2(\register_file[18][30] ),
    .ZN(_07452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12956_ (.A1(_07306_),
    .A2(_07410_),
    .B(_07452_),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12957_ (.A1(_07407_),
    .A2(\register_file[18][31] ),
    .ZN(_07453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12958_ (.A1(_07308_),
    .A2(_07410_),
    .B(_07453_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12959_ (.A1(_06316_),
    .A2(_03854_),
    .ZN(_07454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12960_ (.I(_07454_),
    .Z(_07455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12961_ (.I(_07455_),
    .Z(_07456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12962_ (.I(_07454_),
    .Z(_07457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12963_ (.I(_07457_),
    .Z(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12964_ (.A1(_07458_),
    .A2(\register_file[17][0] ),
    .ZN(_07459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12965_ (.A1(_07230_),
    .A2(_07456_),
    .B(_07459_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12966_ (.A1(_07458_),
    .A2(\register_file[17][1] ),
    .ZN(_07460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12967_ (.A1(_07237_),
    .A2(_07456_),
    .B(_07460_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12968_ (.A1(_07458_),
    .A2(\register_file[17][2] ),
    .ZN(_07461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12969_ (.A1(_07239_),
    .A2(_07456_),
    .B(_07461_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12970_ (.I(_07457_),
    .Z(_07462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12971_ (.A1(_07462_),
    .A2(\register_file[17][3] ),
    .ZN(_07463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12972_ (.A1(_07241_),
    .A2(_07456_),
    .B(_07463_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12973_ (.A1(_07462_),
    .A2(\register_file[17][4] ),
    .ZN(_07464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12974_ (.A1(_07244_),
    .A2(_07456_),
    .B(_07464_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12975_ (.I(_07457_),
    .Z(_07465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12976_ (.I(_07465_),
    .Z(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12977_ (.A1(_07462_),
    .A2(\register_file[17][5] ),
    .ZN(_07467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12978_ (.A1(_07246_),
    .A2(_07466_),
    .B(_07467_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12979_ (.A1(_07462_),
    .A2(\register_file[17][6] ),
    .ZN(_07468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12980_ (.A1(_07250_),
    .A2(_07466_),
    .B(_07468_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12981_ (.A1(_07462_),
    .A2(\register_file[17][7] ),
    .ZN(_07469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12982_ (.A1(_07252_),
    .A2(_07466_),
    .B(_07469_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12983_ (.I(_07457_),
    .Z(_07470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12984_ (.A1(_07470_),
    .A2(\register_file[17][8] ),
    .ZN(_07471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12985_ (.A1(_07254_),
    .A2(_07466_),
    .B(_07471_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12986_ (.A1(_07470_),
    .A2(\register_file[17][9] ),
    .ZN(_07472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12987_ (.A1(_07257_),
    .A2(_07466_),
    .B(_07472_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12988_ (.I(_07465_),
    .Z(_07473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12989_ (.A1(_07470_),
    .A2(\register_file[17][10] ),
    .ZN(_07474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12990_ (.A1(_07259_),
    .A2(_07473_),
    .B(_07474_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12991_ (.A1(_07470_),
    .A2(\register_file[17][11] ),
    .ZN(_07475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12992_ (.A1(_07262_),
    .A2(_07473_),
    .B(_07475_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12993_ (.A1(_07470_),
    .A2(\register_file[17][12] ),
    .ZN(_07476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12994_ (.A1(_07264_),
    .A2(_07473_),
    .B(_07476_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12995_ (.I(_07457_),
    .Z(_07477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12996_ (.A1(_07477_),
    .A2(\register_file[17][13] ),
    .ZN(_07478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12997_ (.A1(_07266_),
    .A2(_07473_),
    .B(_07478_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12998_ (.A1(_07477_),
    .A2(\register_file[17][14] ),
    .ZN(_07479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12999_ (.A1(_07269_),
    .A2(_07473_),
    .B(_07479_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13000_ (.I(_07465_),
    .Z(_07480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13001_ (.A1(_07477_),
    .A2(\register_file[17][15] ),
    .ZN(_07481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13002_ (.A1(_07271_),
    .A2(_07480_),
    .B(_07481_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13003_ (.A1(_07477_),
    .A2(\register_file[17][16] ),
    .ZN(_07482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13004_ (.A1(_07274_),
    .A2(_07480_),
    .B(_07482_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13005_ (.A1(_07477_),
    .A2(\register_file[17][17] ),
    .ZN(_07483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13006_ (.A1(_07276_),
    .A2(_07480_),
    .B(_07483_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13007_ (.I(_07454_),
    .Z(_07484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13008_ (.A1(_07484_),
    .A2(\register_file[17][18] ),
    .ZN(_07485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13009_ (.A1(_07278_),
    .A2(_07480_),
    .B(_07485_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13010_ (.A1(_07484_),
    .A2(\register_file[17][19] ),
    .ZN(_07486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13011_ (.A1(_07281_),
    .A2(_07480_),
    .B(_07486_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13012_ (.I(_07465_),
    .Z(_07487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13013_ (.A1(_07484_),
    .A2(\register_file[17][20] ),
    .ZN(_07488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13014_ (.A1(_07283_),
    .A2(_07487_),
    .B(_07488_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13015_ (.A1(_07484_),
    .A2(\register_file[17][21] ),
    .ZN(_07489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13016_ (.A1(_07286_),
    .A2(_07487_),
    .B(_07489_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13017_ (.A1(_07484_),
    .A2(\register_file[17][22] ),
    .ZN(_07490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13018_ (.A1(_07288_),
    .A2(_07487_),
    .B(_07490_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13019_ (.I(_07454_),
    .Z(_07491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13020_ (.A1(_07491_),
    .A2(\register_file[17][23] ),
    .ZN(_07492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13021_ (.A1(_07290_),
    .A2(_07487_),
    .B(_07492_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13022_ (.A1(_07491_),
    .A2(\register_file[17][24] ),
    .ZN(_07493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13023_ (.A1(_07293_),
    .A2(_07487_),
    .B(_07493_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13024_ (.I(_07465_),
    .Z(_07494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13025_ (.A1(_07491_),
    .A2(\register_file[17][25] ),
    .ZN(_07495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13026_ (.A1(_07295_),
    .A2(_07494_),
    .B(_07495_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13027_ (.A1(_07491_),
    .A2(\register_file[17][26] ),
    .ZN(_07496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13028_ (.A1(_07298_),
    .A2(_07494_),
    .B(_07496_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13029_ (.A1(_07491_),
    .A2(\register_file[17][27] ),
    .ZN(_07497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13030_ (.A1(_07300_),
    .A2(_07494_),
    .B(_07497_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13031_ (.A1(_07455_),
    .A2(\register_file[17][28] ),
    .ZN(_07498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13032_ (.A1(_07302_),
    .A2(_07494_),
    .B(_07498_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13033_ (.A1(_07455_),
    .A2(\register_file[17][29] ),
    .ZN(_07499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13034_ (.A1(_07304_),
    .A2(_07494_),
    .B(_07499_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13035_ (.A1(_07455_),
    .A2(\register_file[17][30] ),
    .ZN(_07500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13036_ (.A1(_07306_),
    .A2(_07458_),
    .B(_07500_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13037_ (.A1(_07455_),
    .A2(\register_file[17][31] ),
    .ZN(_07501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13038_ (.A1(_07308_),
    .A2(_07458_),
    .B(_07501_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13039_ (.I(_06019_),
    .Z(_07502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13040_ (.A1(_06216_),
    .A2(_03854_),
    .ZN(_07503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13041_ (.I(_07503_),
    .Z(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13042_ (.I(_07504_),
    .Z(_07505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13043_ (.I(_07503_),
    .Z(_07506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13044_ (.I(_07506_),
    .Z(_07507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13045_ (.A1(_07507_),
    .A2(\register_file[16][0] ),
    .ZN(_07508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13046_ (.A1(_07502_),
    .A2(_07505_),
    .B(_07508_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13047_ (.I(_06031_),
    .Z(_07509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13048_ (.A1(_07507_),
    .A2(\register_file[16][1] ),
    .ZN(_07510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13049_ (.A1(_07509_),
    .A2(_07505_),
    .B(_07510_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13050_ (.I(_06035_),
    .Z(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13051_ (.A1(_07507_),
    .A2(\register_file[16][2] ),
    .ZN(_07512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13052_ (.A1(_07511_),
    .A2(_07505_),
    .B(_07512_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13053_ (.I(_06039_),
    .Z(_07513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13054_ (.I(_07506_),
    .Z(_07514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13055_ (.A1(_07514_),
    .A2(\register_file[16][3] ),
    .ZN(_07515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13056_ (.A1(_07513_),
    .A2(_07505_),
    .B(_07515_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13057_ (.I(_06044_),
    .Z(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13058_ (.A1(_07514_),
    .A2(\register_file[16][4] ),
    .ZN(_07517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13059_ (.A1(_07516_),
    .A2(_07505_),
    .B(_07517_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13060_ (.I(_06048_),
    .Z(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13061_ (.I(_07506_),
    .Z(_07519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13062_ (.I(_07519_),
    .Z(_07520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13063_ (.A1(_07514_),
    .A2(\register_file[16][5] ),
    .ZN(_07521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13064_ (.A1(_07518_),
    .A2(_07520_),
    .B(_07521_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13065_ (.I(_06054_),
    .Z(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13066_ (.A1(_07514_),
    .A2(\register_file[16][6] ),
    .ZN(_07523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13067_ (.A1(_07522_),
    .A2(_07520_),
    .B(_07523_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13068_ (.I(_06058_),
    .Z(_07524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13069_ (.A1(_07514_),
    .A2(\register_file[16][7] ),
    .ZN(_07525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13070_ (.A1(_07524_),
    .A2(_07520_),
    .B(_07525_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13071_ (.I(_06062_),
    .Z(_07526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13072_ (.I(_07506_),
    .Z(_07527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13073_ (.A1(_07527_),
    .A2(\register_file[16][8] ),
    .ZN(_07528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13074_ (.A1(_07526_),
    .A2(_07520_),
    .B(_07528_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13075_ (.I(_06067_),
    .Z(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13076_ (.A1(_07527_),
    .A2(\register_file[16][9] ),
    .ZN(_07530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13077_ (.A1(_07529_),
    .A2(_07520_),
    .B(_07530_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13078_ (.I(_06071_),
    .Z(_07531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13079_ (.I(_07519_),
    .Z(_07532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13080_ (.A1(_07527_),
    .A2(\register_file[16][10] ),
    .ZN(_07533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13081_ (.A1(_07531_),
    .A2(_07532_),
    .B(_07533_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13082_ (.I(_06076_),
    .Z(_07534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13083_ (.A1(_07527_),
    .A2(\register_file[16][11] ),
    .ZN(_07535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13084_ (.A1(_07534_),
    .A2(_07532_),
    .B(_07535_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13085_ (.I(_06080_),
    .Z(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13086_ (.A1(_07527_),
    .A2(\register_file[16][12] ),
    .ZN(_07537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13087_ (.A1(_07536_),
    .A2(_07532_),
    .B(_07537_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13088_ (.I(_06084_),
    .Z(_07538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13089_ (.I(_07506_),
    .Z(_07539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13090_ (.A1(_07539_),
    .A2(\register_file[16][13] ),
    .ZN(_07540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13091_ (.A1(_07538_),
    .A2(_07532_),
    .B(_07540_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13092_ (.I(_06089_),
    .Z(_07541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13093_ (.A1(_07539_),
    .A2(\register_file[16][14] ),
    .ZN(_07542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13094_ (.A1(_07541_),
    .A2(_07532_),
    .B(_07542_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13095_ (.I(_06093_),
    .Z(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13096_ (.I(_07519_),
    .Z(_07544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13097_ (.A1(_07539_),
    .A2(\register_file[16][15] ),
    .ZN(_07545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13098_ (.A1(_07543_),
    .A2(_07544_),
    .B(_07545_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13099_ (.I(_06098_),
    .Z(_07546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13100_ (.A1(_07539_),
    .A2(\register_file[16][16] ),
    .ZN(_07547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13101_ (.A1(_07546_),
    .A2(_07544_),
    .B(_07547_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13102_ (.I(_06102_),
    .Z(_07548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13103_ (.A1(_07539_),
    .A2(\register_file[16][17] ),
    .ZN(_07549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13104_ (.A1(_07548_),
    .A2(_07544_),
    .B(_07549_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13105_ (.I(_06106_),
    .Z(_07550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13106_ (.I(_07503_),
    .Z(_07551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13107_ (.A1(_07551_),
    .A2(\register_file[16][18] ),
    .ZN(_07552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13108_ (.A1(_07550_),
    .A2(_07544_),
    .B(_07552_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13109_ (.I(_06111_),
    .Z(_07553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13110_ (.A1(_07551_),
    .A2(\register_file[16][19] ),
    .ZN(_07554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13111_ (.A1(_07553_),
    .A2(_07544_),
    .B(_07554_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13112_ (.I(_06115_),
    .Z(_07555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13113_ (.I(_07519_),
    .Z(_07556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13114_ (.A1(_07551_),
    .A2(\register_file[16][20] ),
    .ZN(_07557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13115_ (.A1(_07555_),
    .A2(_07556_),
    .B(_07557_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13116_ (.I(_06120_),
    .Z(_07558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13117_ (.A1(_07551_),
    .A2(\register_file[16][21] ),
    .ZN(_07559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13118_ (.A1(_07558_),
    .A2(_07556_),
    .B(_07559_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13119_ (.I(_06124_),
    .Z(_07560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13120_ (.A1(_07551_),
    .A2(\register_file[16][22] ),
    .ZN(_07561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13121_ (.A1(_07560_),
    .A2(_07556_),
    .B(_07561_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13122_ (.I(_06128_),
    .Z(_07562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13123_ (.I(_07503_),
    .Z(_07563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13124_ (.A1(_07563_),
    .A2(\register_file[16][23] ),
    .ZN(_07564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13125_ (.A1(_07562_),
    .A2(_07556_),
    .B(_07564_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13126_ (.I(_06133_),
    .Z(_07565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13127_ (.A1(_07563_),
    .A2(\register_file[16][24] ),
    .ZN(_07566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13128_ (.A1(_07565_),
    .A2(_07556_),
    .B(_07566_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13129_ (.I(_06137_),
    .Z(_07567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13130_ (.I(_07519_),
    .Z(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13131_ (.A1(_07563_),
    .A2(\register_file[16][25] ),
    .ZN(_07569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13132_ (.A1(_07567_),
    .A2(_07568_),
    .B(_07569_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13133_ (.I(_06142_),
    .Z(_07570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13134_ (.A1(_07563_),
    .A2(\register_file[16][26] ),
    .ZN(_07571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13135_ (.A1(_07570_),
    .A2(_07568_),
    .B(_07571_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13136_ (.I(_06146_),
    .Z(_07572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13137_ (.A1(_07563_),
    .A2(\register_file[16][27] ),
    .ZN(_07573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13138_ (.A1(_07572_),
    .A2(_07568_),
    .B(_07573_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13139_ (.I(_06150_),
    .Z(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13140_ (.A1(_07504_),
    .A2(\register_file[16][28] ),
    .ZN(_07575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13141_ (.A1(_07574_),
    .A2(_07568_),
    .B(_07575_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13142_ (.I(_06154_),
    .Z(_07576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13143_ (.A1(_07504_),
    .A2(\register_file[16][29] ),
    .ZN(_07577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13144_ (.A1(_07576_),
    .A2(_07568_),
    .B(_07577_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13145_ (.I(_06158_),
    .Z(_07578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13146_ (.A1(_07504_),
    .A2(\register_file[16][30] ),
    .ZN(_07579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13147_ (.A1(_07578_),
    .A2(_07507_),
    .B(_07579_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13148_ (.I(_06162_),
    .Z(_07580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13149_ (.A1(_07504_),
    .A2(\register_file[16][31] ),
    .ZN(_07581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13150_ (.A1(_07580_),
    .A2(_07507_),
    .B(_07581_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13151_ (.A1(_06265_),
    .A2(_03875_),
    .ZN(_07582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13152_ (.I(_07582_),
    .Z(_07583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13153_ (.I(_07583_),
    .Z(_07584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13154_ (.I(_07582_),
    .Z(_07585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13155_ (.I(_07585_),
    .Z(_07586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13156_ (.A1(_07586_),
    .A2(\register_file[15][0] ),
    .ZN(_07587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13157_ (.A1(_07502_),
    .A2(_07584_),
    .B(_07587_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13158_ (.A1(_07586_),
    .A2(\register_file[15][1] ),
    .ZN(_07588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13159_ (.A1(_07509_),
    .A2(_07584_),
    .B(_07588_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13160_ (.A1(_07586_),
    .A2(\register_file[15][2] ),
    .ZN(_07589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13161_ (.A1(_07511_),
    .A2(_07584_),
    .B(_07589_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13162_ (.I(_07585_),
    .Z(_07590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13163_ (.A1(_07590_),
    .A2(\register_file[15][3] ),
    .ZN(_07591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13164_ (.A1(_07513_),
    .A2(_07584_),
    .B(_07591_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13165_ (.A1(_07590_),
    .A2(\register_file[15][4] ),
    .ZN(_07592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13166_ (.A1(_07516_),
    .A2(_07584_),
    .B(_07592_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13167_ (.I(_07585_),
    .Z(_07593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13168_ (.I(_07593_),
    .Z(_07594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13169_ (.A1(_07590_),
    .A2(\register_file[15][5] ),
    .ZN(_07595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13170_ (.A1(_07518_),
    .A2(_07594_),
    .B(_07595_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13171_ (.A1(_07590_),
    .A2(\register_file[15][6] ),
    .ZN(_07596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13172_ (.A1(_07522_),
    .A2(_07594_),
    .B(_07596_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13173_ (.A1(_07590_),
    .A2(\register_file[15][7] ),
    .ZN(_07597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13174_ (.A1(_07524_),
    .A2(_07594_),
    .B(_07597_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13175_ (.I(_07585_),
    .Z(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13176_ (.A1(_07598_),
    .A2(\register_file[15][8] ),
    .ZN(_07599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13177_ (.A1(_07526_),
    .A2(_07594_),
    .B(_07599_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13178_ (.A1(_07598_),
    .A2(\register_file[15][9] ),
    .ZN(_07600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13179_ (.A1(_07529_),
    .A2(_07594_),
    .B(_07600_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13180_ (.I(_07593_),
    .Z(_07601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13181_ (.A1(_07598_),
    .A2(\register_file[15][10] ),
    .ZN(_07602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13182_ (.A1(_07531_),
    .A2(_07601_),
    .B(_07602_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13183_ (.A1(_07598_),
    .A2(\register_file[15][11] ),
    .ZN(_07603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13184_ (.A1(_07534_),
    .A2(_07601_),
    .B(_07603_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13185_ (.A1(_07598_),
    .A2(\register_file[15][12] ),
    .ZN(_07604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13186_ (.A1(_07536_),
    .A2(_07601_),
    .B(_07604_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13187_ (.I(_07585_),
    .Z(_07605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13188_ (.A1(_07605_),
    .A2(\register_file[15][13] ),
    .ZN(_07606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13189_ (.A1(_07538_),
    .A2(_07601_),
    .B(_07606_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13190_ (.A1(_07605_),
    .A2(\register_file[15][14] ),
    .ZN(_07607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13191_ (.A1(_07541_),
    .A2(_07601_),
    .B(_07607_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13192_ (.I(_07593_),
    .Z(_07608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13193_ (.A1(_07605_),
    .A2(\register_file[15][15] ),
    .ZN(_07609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13194_ (.A1(_07543_),
    .A2(_07608_),
    .B(_07609_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13195_ (.A1(_07605_),
    .A2(\register_file[15][16] ),
    .ZN(_07610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13196_ (.A1(_07546_),
    .A2(_07608_),
    .B(_07610_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13197_ (.A1(_07605_),
    .A2(\register_file[15][17] ),
    .ZN(_07611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13198_ (.A1(_07548_),
    .A2(_07608_),
    .B(_07611_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13199_ (.I(_07582_),
    .Z(_07612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13200_ (.A1(_07612_),
    .A2(\register_file[15][18] ),
    .ZN(_07613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13201_ (.A1(_07550_),
    .A2(_07608_),
    .B(_07613_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13202_ (.A1(_07612_),
    .A2(\register_file[15][19] ),
    .ZN(_07614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13203_ (.A1(_07553_),
    .A2(_07608_),
    .B(_07614_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13204_ (.I(_07593_),
    .Z(_07615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13205_ (.A1(_07612_),
    .A2(\register_file[15][20] ),
    .ZN(_07616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13206_ (.A1(_07555_),
    .A2(_07615_),
    .B(_07616_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13207_ (.A1(_07612_),
    .A2(\register_file[15][21] ),
    .ZN(_07617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13208_ (.A1(_07558_),
    .A2(_07615_),
    .B(_07617_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13209_ (.A1(_07612_),
    .A2(\register_file[15][22] ),
    .ZN(_07618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13210_ (.A1(_07560_),
    .A2(_07615_),
    .B(_07618_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13211_ (.I(_07582_),
    .Z(_07619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13212_ (.A1(_07619_),
    .A2(\register_file[15][23] ),
    .ZN(_07620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13213_ (.A1(_07562_),
    .A2(_07615_),
    .B(_07620_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13214_ (.A1(_07619_),
    .A2(\register_file[15][24] ),
    .ZN(_07621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13215_ (.A1(_07565_),
    .A2(_07615_),
    .B(_07621_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13216_ (.I(_07593_),
    .Z(_07622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13217_ (.A1(_07619_),
    .A2(\register_file[15][25] ),
    .ZN(_07623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13218_ (.A1(_07567_),
    .A2(_07622_),
    .B(_07623_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13219_ (.A1(_07619_),
    .A2(\register_file[15][26] ),
    .ZN(_07624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13220_ (.A1(_07570_),
    .A2(_07622_),
    .B(_07624_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13221_ (.A1(_07619_),
    .A2(\register_file[15][27] ),
    .ZN(_07625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13222_ (.A1(_07572_),
    .A2(_07622_),
    .B(_07625_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13223_ (.A1(_07583_),
    .A2(\register_file[15][28] ),
    .ZN(_07626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13224_ (.A1(_07574_),
    .A2(_07622_),
    .B(_07626_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13225_ (.A1(_07583_),
    .A2(\register_file[15][29] ),
    .ZN(_07627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13226_ (.A1(_07576_),
    .A2(_07622_),
    .B(_07627_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13227_ (.A1(_07583_),
    .A2(\register_file[15][30] ),
    .ZN(_07628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13228_ (.A1(_07578_),
    .A2(_07586_),
    .B(_07628_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13229_ (.A1(_07583_),
    .A2(\register_file[15][31] ),
    .ZN(_07629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13230_ (.A1(_07580_),
    .A2(_07586_),
    .B(_07629_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13231_ (.A1(_06023_),
    .A2(_03875_),
    .ZN(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13232_ (.I(_07630_),
    .Z(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13233_ (.I(_07631_),
    .Z(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13234_ (.I(_07630_),
    .Z(_07633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13235_ (.I(_07633_),
    .Z(_07634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13236_ (.A1(_07634_),
    .A2(\register_file[14][0] ),
    .ZN(_07635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13237_ (.A1(_07502_),
    .A2(_07632_),
    .B(_07635_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13238_ (.A1(_07634_),
    .A2(\register_file[14][1] ),
    .ZN(_07636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13239_ (.A1(_07509_),
    .A2(_07632_),
    .B(_07636_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13240_ (.A1(_07634_),
    .A2(\register_file[14][2] ),
    .ZN(_07637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13241_ (.A1(_07511_),
    .A2(_07632_),
    .B(_07637_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13242_ (.I(_07633_),
    .Z(_07638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13243_ (.A1(_07638_),
    .A2(\register_file[14][3] ),
    .ZN(_07639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13244_ (.A1(_07513_),
    .A2(_07632_),
    .B(_07639_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13245_ (.A1(_07638_),
    .A2(\register_file[14][4] ),
    .ZN(_07640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13246_ (.A1(_07516_),
    .A2(_07632_),
    .B(_07640_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13247_ (.I(_07633_),
    .Z(_07641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13248_ (.I(_07641_),
    .Z(_07642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13249_ (.A1(_07638_),
    .A2(\register_file[14][5] ),
    .ZN(_07643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13250_ (.A1(_07518_),
    .A2(_07642_),
    .B(_07643_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13251_ (.A1(_07638_),
    .A2(\register_file[14][6] ),
    .ZN(_07644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13252_ (.A1(_07522_),
    .A2(_07642_),
    .B(_07644_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13253_ (.A1(_07638_),
    .A2(\register_file[14][7] ),
    .ZN(_07645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13254_ (.A1(_07524_),
    .A2(_07642_),
    .B(_07645_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13255_ (.I(_07633_),
    .Z(_07646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13256_ (.A1(_07646_),
    .A2(\register_file[14][8] ),
    .ZN(_07647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13257_ (.A1(_07526_),
    .A2(_07642_),
    .B(_07647_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13258_ (.A1(_07646_),
    .A2(\register_file[14][9] ),
    .ZN(_07648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13259_ (.A1(_07529_),
    .A2(_07642_),
    .B(_07648_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13260_ (.I(_07641_),
    .Z(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13261_ (.A1(_07646_),
    .A2(\register_file[14][10] ),
    .ZN(_07650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13262_ (.A1(_07531_),
    .A2(_07649_),
    .B(_07650_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13263_ (.A1(_07646_),
    .A2(\register_file[14][11] ),
    .ZN(_07651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13264_ (.A1(_07534_),
    .A2(_07649_),
    .B(_07651_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13265_ (.A1(_07646_),
    .A2(\register_file[14][12] ),
    .ZN(_07652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13266_ (.A1(_07536_),
    .A2(_07649_),
    .B(_07652_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13267_ (.I(_07633_),
    .Z(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13268_ (.A1(_07653_),
    .A2(\register_file[14][13] ),
    .ZN(_07654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13269_ (.A1(_07538_),
    .A2(_07649_),
    .B(_07654_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13270_ (.A1(_07653_),
    .A2(\register_file[14][14] ),
    .ZN(_07655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13271_ (.A1(_07541_),
    .A2(_07649_),
    .B(_07655_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13272_ (.I(_07641_),
    .Z(_07656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13273_ (.A1(_07653_),
    .A2(\register_file[14][15] ),
    .ZN(_07657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13274_ (.A1(_07543_),
    .A2(_07656_),
    .B(_07657_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13275_ (.A1(_07653_),
    .A2(\register_file[14][16] ),
    .ZN(_07658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13276_ (.A1(_07546_),
    .A2(_07656_),
    .B(_07658_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13277_ (.A1(_07653_),
    .A2(\register_file[14][17] ),
    .ZN(_07659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13278_ (.A1(_07548_),
    .A2(_07656_),
    .B(_07659_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13279_ (.I(_07630_),
    .Z(_07660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13280_ (.A1(_07660_),
    .A2(\register_file[14][18] ),
    .ZN(_07661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13281_ (.A1(_07550_),
    .A2(_07656_),
    .B(_07661_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13282_ (.A1(_07660_),
    .A2(\register_file[14][19] ),
    .ZN(_07662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13283_ (.A1(_07553_),
    .A2(_07656_),
    .B(_07662_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13284_ (.I(_07641_),
    .Z(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13285_ (.A1(_07660_),
    .A2(\register_file[14][20] ),
    .ZN(_07664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13286_ (.A1(_07555_),
    .A2(_07663_),
    .B(_07664_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13287_ (.A1(_07660_),
    .A2(\register_file[14][21] ),
    .ZN(_07665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13288_ (.A1(_07558_),
    .A2(_07663_),
    .B(_07665_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13289_ (.A1(_07660_),
    .A2(\register_file[14][22] ),
    .ZN(_07666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13290_ (.A1(_07560_),
    .A2(_07663_),
    .B(_07666_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13291_ (.I(_07630_),
    .Z(_07667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13292_ (.A1(_07667_),
    .A2(\register_file[14][23] ),
    .ZN(_07668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13293_ (.A1(_07562_),
    .A2(_07663_),
    .B(_07668_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13294_ (.A1(_07667_),
    .A2(\register_file[14][24] ),
    .ZN(_07669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13295_ (.A1(_07565_),
    .A2(_07663_),
    .B(_07669_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13296_ (.I(_07641_),
    .Z(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13297_ (.A1(_07667_),
    .A2(\register_file[14][25] ),
    .ZN(_07671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13298_ (.A1(_07567_),
    .A2(_07670_),
    .B(_07671_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13299_ (.A1(_07667_),
    .A2(\register_file[14][26] ),
    .ZN(_07672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13300_ (.A1(_07570_),
    .A2(_07670_),
    .B(_07672_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13301_ (.A1(_07667_),
    .A2(\register_file[14][27] ),
    .ZN(_07673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13302_ (.A1(_07572_),
    .A2(_07670_),
    .B(_07673_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13303_ (.A1(_07631_),
    .A2(\register_file[14][28] ),
    .ZN(_07674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13304_ (.A1(_07574_),
    .A2(_07670_),
    .B(_07674_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13305_ (.A1(_07631_),
    .A2(\register_file[14][29] ),
    .ZN(_07675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13306_ (.A1(_07576_),
    .A2(_07670_),
    .B(_07675_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13307_ (.A1(_07631_),
    .A2(\register_file[14][30] ),
    .ZN(_07676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13308_ (.A1(_07578_),
    .A2(_07634_),
    .B(_07676_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13309_ (.A1(_07631_),
    .A2(\register_file[14][31] ),
    .ZN(_07677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13310_ (.A1(_07580_),
    .A2(_07634_),
    .B(_07677_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13311_ (.A1(_06316_),
    .A2(_03815_),
    .ZN(_07678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13312_ (.I(_07678_),
    .Z(_07679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13313_ (.I(_07679_),
    .Z(_07680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13314_ (.I(_07678_),
    .Z(_07681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13315_ (.I(_07681_),
    .Z(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13316_ (.A1(_07682_),
    .A2(\register_file[29][0] ),
    .ZN(_07683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13317_ (.A1(_07502_),
    .A2(_07680_),
    .B(_07683_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13318_ (.A1(_07682_),
    .A2(\register_file[29][1] ),
    .ZN(_07684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13319_ (.A1(_07509_),
    .A2(_07680_),
    .B(_07684_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13320_ (.A1(_07682_),
    .A2(\register_file[29][2] ),
    .ZN(_07685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13321_ (.A1(_07511_),
    .A2(_07680_),
    .B(_07685_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13322_ (.I(_07681_),
    .Z(_07686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13323_ (.A1(_07686_),
    .A2(\register_file[29][3] ),
    .ZN(_07687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13324_ (.A1(_07513_),
    .A2(_07680_),
    .B(_07687_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13325_ (.A1(_07686_),
    .A2(\register_file[29][4] ),
    .ZN(_07688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13326_ (.A1(_07516_),
    .A2(_07680_),
    .B(_07688_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13327_ (.I(_07681_),
    .Z(_07689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13328_ (.I(_07689_),
    .Z(_07690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13329_ (.A1(_07686_),
    .A2(\register_file[29][5] ),
    .ZN(_07691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13330_ (.A1(_07518_),
    .A2(_07690_),
    .B(_07691_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13331_ (.A1(_07686_),
    .A2(\register_file[29][6] ),
    .ZN(_07692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13332_ (.A1(_07522_),
    .A2(_07690_),
    .B(_07692_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13333_ (.A1(_07686_),
    .A2(\register_file[29][7] ),
    .ZN(_07693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13334_ (.A1(_07524_),
    .A2(_07690_),
    .B(_07693_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13335_ (.I(_07681_),
    .Z(_07694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13336_ (.A1(_07694_),
    .A2(\register_file[29][8] ),
    .ZN(_07695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13337_ (.A1(_07526_),
    .A2(_07690_),
    .B(_07695_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13338_ (.A1(_07694_),
    .A2(\register_file[29][9] ),
    .ZN(_07696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13339_ (.A1(_07529_),
    .A2(_07690_),
    .B(_07696_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13340_ (.I(_07689_),
    .Z(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13341_ (.A1(_07694_),
    .A2(\register_file[29][10] ),
    .ZN(_07698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13342_ (.A1(_07531_),
    .A2(_07697_),
    .B(_07698_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13343_ (.A1(_07694_),
    .A2(\register_file[29][11] ),
    .ZN(_07699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13344_ (.A1(_07534_),
    .A2(_07697_),
    .B(_07699_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13345_ (.A1(_07694_),
    .A2(\register_file[29][12] ),
    .ZN(_07700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13346_ (.A1(_07536_),
    .A2(_07697_),
    .B(_07700_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13347_ (.I(_07681_),
    .Z(_07701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13348_ (.A1(_07701_),
    .A2(\register_file[29][13] ),
    .ZN(_07702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13349_ (.A1(_07538_),
    .A2(_07697_),
    .B(_07702_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13350_ (.A1(_07701_),
    .A2(\register_file[29][14] ),
    .ZN(_07703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13351_ (.A1(_07541_),
    .A2(_07697_),
    .B(_07703_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13352_ (.I(_07689_),
    .Z(_07704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13353_ (.A1(_07701_),
    .A2(\register_file[29][15] ),
    .ZN(_07705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13354_ (.A1(_07543_),
    .A2(_07704_),
    .B(_07705_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13355_ (.A1(_07701_),
    .A2(\register_file[29][16] ),
    .ZN(_07706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13356_ (.A1(_07546_),
    .A2(_07704_),
    .B(_07706_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13357_ (.A1(_07701_),
    .A2(\register_file[29][17] ),
    .ZN(_07707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13358_ (.A1(_07548_),
    .A2(_07704_),
    .B(_07707_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13359_ (.I(_07678_),
    .Z(_07708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13360_ (.A1(_07708_),
    .A2(\register_file[29][18] ),
    .ZN(_07709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13361_ (.A1(_07550_),
    .A2(_07704_),
    .B(_07709_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13362_ (.A1(_07708_),
    .A2(\register_file[29][19] ),
    .ZN(_07710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13363_ (.A1(_07553_),
    .A2(_07704_),
    .B(_07710_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13364_ (.I(_07689_),
    .Z(_07711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13365_ (.A1(_07708_),
    .A2(\register_file[29][20] ),
    .ZN(_07712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13366_ (.A1(_07555_),
    .A2(_07711_),
    .B(_07712_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13367_ (.A1(_07708_),
    .A2(\register_file[29][21] ),
    .ZN(_07713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13368_ (.A1(_07558_),
    .A2(_07711_),
    .B(_07713_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13369_ (.A1(_07708_),
    .A2(\register_file[29][22] ),
    .ZN(_07714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13370_ (.A1(_07560_),
    .A2(_07711_),
    .B(_07714_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13371_ (.I(_07678_),
    .Z(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13372_ (.A1(_07715_),
    .A2(\register_file[29][23] ),
    .ZN(_07716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13373_ (.A1(_07562_),
    .A2(_07711_),
    .B(_07716_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13374_ (.A1(_07715_),
    .A2(\register_file[29][24] ),
    .ZN(_07717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13375_ (.A1(_07565_),
    .A2(_07711_),
    .B(_07717_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13376_ (.I(_07689_),
    .Z(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13377_ (.A1(_07715_),
    .A2(\register_file[29][25] ),
    .ZN(_07719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13378_ (.A1(_07567_),
    .A2(_07718_),
    .B(_07719_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13379_ (.A1(_07715_),
    .A2(\register_file[29][26] ),
    .ZN(_07720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13380_ (.A1(_07570_),
    .A2(_07718_),
    .B(_07720_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13381_ (.A1(_07715_),
    .A2(\register_file[29][27] ),
    .ZN(_07721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13382_ (.A1(_07572_),
    .A2(_07718_),
    .B(_07721_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13383_ (.A1(_07679_),
    .A2(\register_file[29][28] ),
    .ZN(_07722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13384_ (.A1(_07574_),
    .A2(_07718_),
    .B(_07722_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13385_ (.A1(_07679_),
    .A2(\register_file[29][29] ),
    .ZN(_07723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13386_ (.A1(_07576_),
    .A2(_07718_),
    .B(_07723_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13387_ (.A1(_07679_),
    .A2(\register_file[29][30] ),
    .ZN(_07724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13388_ (.A1(_07578_),
    .A2(_07682_),
    .B(_07724_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13389_ (.A1(_07679_),
    .A2(\register_file[29][31] ),
    .ZN(_07725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13390_ (.A1(_07580_),
    .A2(_07682_),
    .B(_07725_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13391_ (.A1(_06316_),
    .A2(_03893_),
    .ZN(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13392_ (.I(_07726_),
    .Z(_07727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13393_ (.I(_07727_),
    .Z(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13394_ (.I(_07726_),
    .Z(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13395_ (.I(_07729_),
    .Z(_07730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13396_ (.A1(_07730_),
    .A2(\register_file[9][0] ),
    .ZN(_07731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13397_ (.A1(_07502_),
    .A2(_07728_),
    .B(_07731_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13398_ (.A1(_07730_),
    .A2(\register_file[9][1] ),
    .ZN(_07732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13399_ (.A1(_07509_),
    .A2(_07728_),
    .B(_07732_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13400_ (.A1(_07730_),
    .A2(\register_file[9][2] ),
    .ZN(_07733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13401_ (.A1(_07511_),
    .A2(_07728_),
    .B(_07733_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13402_ (.I(_07729_),
    .Z(_07734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13403_ (.A1(_07734_),
    .A2(\register_file[9][3] ),
    .ZN(_07735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13404_ (.A1(_07513_),
    .A2(_07728_),
    .B(_07735_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13405_ (.A1(_07734_),
    .A2(\register_file[9][4] ),
    .ZN(_07736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13406_ (.A1(_07516_),
    .A2(_07728_),
    .B(_07736_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13407_ (.I(_07729_),
    .Z(_07737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13408_ (.I(_07737_),
    .Z(_07738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13409_ (.A1(_07734_),
    .A2(\register_file[9][5] ),
    .ZN(_07739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13410_ (.A1(_07518_),
    .A2(_07738_),
    .B(_07739_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13411_ (.A1(_07734_),
    .A2(\register_file[9][6] ),
    .ZN(_07740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13412_ (.A1(_07522_),
    .A2(_07738_),
    .B(_07740_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13413_ (.A1(_07734_),
    .A2(\register_file[9][7] ),
    .ZN(_07741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13414_ (.A1(_07524_),
    .A2(_07738_),
    .B(_07741_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13415_ (.I(_07729_),
    .Z(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13416_ (.A1(_07742_),
    .A2(\register_file[9][8] ),
    .ZN(_07743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13417_ (.A1(_07526_),
    .A2(_07738_),
    .B(_07743_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13418_ (.A1(_07742_),
    .A2(\register_file[9][9] ),
    .ZN(_07744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13419_ (.A1(_07529_),
    .A2(_07738_),
    .B(_07744_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13420_ (.I(_07737_),
    .Z(_07745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13421_ (.A1(_07742_),
    .A2(\register_file[9][10] ),
    .ZN(_07746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13422_ (.A1(_07531_),
    .A2(_07745_),
    .B(_07746_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13423_ (.A1(_07742_),
    .A2(\register_file[9][11] ),
    .ZN(_07747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13424_ (.A1(_07534_),
    .A2(_07745_),
    .B(_07747_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13425_ (.A1(_07742_),
    .A2(\register_file[9][12] ),
    .ZN(_07748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13426_ (.A1(_07536_),
    .A2(_07745_),
    .B(_07748_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13427_ (.I(_07729_),
    .Z(_07749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13428_ (.A1(_07749_),
    .A2(\register_file[9][13] ),
    .ZN(_07750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13429_ (.A1(_07538_),
    .A2(_07745_),
    .B(_07750_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13430_ (.A1(_07749_),
    .A2(\register_file[9][14] ),
    .ZN(_07751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13431_ (.A1(_07541_),
    .A2(_07745_),
    .B(_07751_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13432_ (.I(_07737_),
    .Z(_07752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13433_ (.A1(_07749_),
    .A2(\register_file[9][15] ),
    .ZN(_07753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13434_ (.A1(_07543_),
    .A2(_07752_),
    .B(_07753_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13435_ (.A1(_07749_),
    .A2(\register_file[9][16] ),
    .ZN(_07754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13436_ (.A1(_07546_),
    .A2(_07752_),
    .B(_07754_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13437_ (.A1(_07749_),
    .A2(\register_file[9][17] ),
    .ZN(_07755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13438_ (.A1(_07548_),
    .A2(_07752_),
    .B(_07755_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13439_ (.I(_07726_),
    .Z(_07756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13440_ (.A1(_07756_),
    .A2(\register_file[9][18] ),
    .ZN(_07757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13441_ (.A1(_07550_),
    .A2(_07752_),
    .B(_07757_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13442_ (.A1(_07756_),
    .A2(\register_file[9][19] ),
    .ZN(_07758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13443_ (.A1(_07553_),
    .A2(_07752_),
    .B(_07758_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13444_ (.I(_07737_),
    .Z(_07759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13445_ (.A1(_07756_),
    .A2(\register_file[9][20] ),
    .ZN(_07760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13446_ (.A1(_07555_),
    .A2(_07759_),
    .B(_07760_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13447_ (.A1(_07756_),
    .A2(\register_file[9][21] ),
    .ZN(_07761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13448_ (.A1(_07558_),
    .A2(_07759_),
    .B(_07761_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13449_ (.A1(_07756_),
    .A2(\register_file[9][22] ),
    .ZN(_07762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13450_ (.A1(_07560_),
    .A2(_07759_),
    .B(_07762_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13451_ (.I(_07726_),
    .Z(_07763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13452_ (.A1(_07763_),
    .A2(\register_file[9][23] ),
    .ZN(_07764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13453_ (.A1(_07562_),
    .A2(_07759_),
    .B(_07764_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13454_ (.A1(_07763_),
    .A2(\register_file[9][24] ),
    .ZN(_07765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13455_ (.A1(_07565_),
    .A2(_07759_),
    .B(_07765_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13456_ (.I(_07737_),
    .Z(_07766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13457_ (.A1(_07763_),
    .A2(\register_file[9][25] ),
    .ZN(_07767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13458_ (.A1(_07567_),
    .A2(_07766_),
    .B(_07767_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13459_ (.A1(_07763_),
    .A2(\register_file[9][26] ),
    .ZN(_07768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13460_ (.A1(_07570_),
    .A2(_07766_),
    .B(_07768_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13461_ (.A1(_07763_),
    .A2(\register_file[9][27] ),
    .ZN(_07769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13462_ (.A1(_07572_),
    .A2(_07766_),
    .B(_07769_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13463_ (.A1(_07727_),
    .A2(\register_file[9][28] ),
    .ZN(_07770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13464_ (.A1(_07574_),
    .A2(_07766_),
    .B(_07770_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13465_ (.A1(_07727_),
    .A2(\register_file[9][29] ),
    .ZN(_07771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13466_ (.A1(_07576_),
    .A2(_07766_),
    .B(_07771_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13467_ (.A1(_07727_),
    .A2(\register_file[9][30] ),
    .ZN(_07772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13468_ (.A1(_07578_),
    .A2(_07730_),
    .B(_07772_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13469_ (.A1(_07727_),
    .A2(\register_file[9][31] ),
    .ZN(_07773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13470_ (.A1(_07580_),
    .A2(_07730_),
    .B(_07773_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13471_ (.I(net6),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13472_ (.I(_00992_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13473_ (.I(_00993_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13474_ (.I(_00994_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13475_ (.A1(_00995_),
    .A2(\register_file[16][0] ),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _13476_ (.I(net6),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _13477_ (.I(_00997_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _13478_ (.I(_00998_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13479_ (.I(_00999_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13480_ (.A1(_01000_),
    .A2(\register_file[17][0] ),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13481_ (.A1(_00996_),
    .A2(_01001_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13482_ (.A1(net7),
    .A2(net8),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13483_ (.I(_01003_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13484_ (.I(_01004_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13485_ (.I(_01005_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13486_ (.A1(_01002_),
    .A2(_01006_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13487_ (.I(net9),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13488_ (.I(_01008_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13489_ (.I(_01009_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13490_ (.I(_01010_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13491_ (.A1(_01007_),
    .A2(_01011_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _13492_ (.I(_00997_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13493_ (.I(_01013_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13494_ (.I(_01014_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13495_ (.A1(_01015_),
    .A2(\register_file[19][0] ),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13496_ (.I(_00992_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13497_ (.I(_01017_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13498_ (.I(_01018_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13499_ (.A1(_01019_),
    .A2(\register_file[18][0] ),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13500_ (.I(net8),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _13501_ (.I(_01021_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13502_ (.I(net7),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13503_ (.A1(_01022_),
    .A2(_01023_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13504_ (.I(_01024_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13505_ (.I(_01025_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13506_ (.A1(_01016_),
    .A2(_01020_),
    .B(_01026_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13507_ (.A1(_01012_),
    .A2(_01027_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13508_ (.I(_00992_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13509_ (.I(_01029_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13510_ (.I(_01030_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13511_ (.A1(_01031_),
    .A2(\register_file[20][0] ),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13512_ (.I(_01023_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13513_ (.I(_01033_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13514_ (.I(_01034_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13515_ (.I(_01035_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13516_ (.I(_00997_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13517_ (.I(_01037_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13518_ (.I(_01038_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13519_ (.A1(_01039_),
    .A2(\register_file[21][0] ),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13520_ (.A1(_01032_),
    .A2(_01036_),
    .A3(_01040_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13521_ (.I(_01017_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13522_ (.I(_01042_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13523_ (.A1(_01043_),
    .A2(\register_file[22][0] ),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13524_ (.I(_01023_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13525_ (.I(_01045_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13526_ (.I(_01037_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13527_ (.I(_01047_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13528_ (.A1(_01048_),
    .A2(\register_file[23][0] ),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13529_ (.A1(_01044_),
    .A2(_01046_),
    .A3(_01049_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13530_ (.I(_01021_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13531_ (.I(_01051_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13532_ (.A1(_01041_),
    .A2(_01050_),
    .A3(_01052_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13533_ (.A1(_01028_),
    .A2(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13534_ (.I(_00993_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13535_ (.I(_01055_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13536_ (.A1(_01056_),
    .A2(\register_file[24][0] ),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13537_ (.I(_00998_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13538_ (.I(_01058_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13539_ (.A1(_01059_),
    .A2(\register_file[25][0] ),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13540_ (.A1(_01057_),
    .A2(_01060_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13541_ (.I(_01004_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13542_ (.I(_01062_),
    .Z(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13543_ (.A1(_01061_),
    .A2(_01063_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13544_ (.I(net9),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13545_ (.I(_01065_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13546_ (.A1(_01064_),
    .A2(_01066_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13547_ (.I(_01013_),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13548_ (.I(_01068_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13549_ (.A1(_01069_),
    .A2(\register_file[27][0] ),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13550_ (.I(_01017_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13551_ (.I(_01071_),
    .Z(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13552_ (.A1(_01072_),
    .A2(\register_file[26][0] ),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13553_ (.I(_01024_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13554_ (.I(_01074_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13555_ (.I(_01075_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13556_ (.A1(_01070_),
    .A2(_01073_),
    .B(_01076_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13557_ (.A1(_01067_),
    .A2(_01077_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13558_ (.I(_00992_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13559_ (.I(_01079_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13560_ (.I(_01080_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13561_ (.A1(_01081_),
    .A2(\register_file[28][0] ),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13562_ (.I(_01034_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13563_ (.I(_01083_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13564_ (.I(_01037_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13565_ (.I(_01085_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13566_ (.A1(_01086_),
    .A2(\register_file[29][0] ),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13567_ (.A1(_01082_),
    .A2(_01084_),
    .A3(_01087_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13568_ (.I(_01029_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13569_ (.I(_01089_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13570_ (.A1(_01090_),
    .A2(\register_file[30][0] ),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13571_ (.I(_01023_),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13572_ (.I(_01092_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13573_ (.I(_01093_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13574_ (.I(_00997_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13575_ (.I(_01095_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13576_ (.I(_01096_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13577_ (.A1(_01097_),
    .A2(\register_file[31][0] ),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13578_ (.A1(_01091_),
    .A2(_01094_),
    .A3(_01098_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13579_ (.I(_01051_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13580_ (.I(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13581_ (.A1(_01088_),
    .A2(_01099_),
    .A3(_01101_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13582_ (.A1(_01078_),
    .A2(_01102_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13583_ (.I(net10),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13584_ (.I(_01104_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13585_ (.A1(_01054_),
    .A2(_01103_),
    .A3(_01105_),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13586_ (.I(_00993_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13587_ (.I(_01107_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13588_ (.A1(_01108_),
    .A2(\register_file[8][0] ),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13589_ (.I(_00997_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13590_ (.I(_01110_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13591_ (.A1(_01111_),
    .A2(\register_file[9][0] ),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13592_ (.A1(_01109_),
    .A2(_01112_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13593_ (.I(_01004_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13594_ (.I(_01114_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13595_ (.A1(_01113_),
    .A2(_01115_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13596_ (.I(_01065_),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13597_ (.A1(_01116_),
    .A2(_01117_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13598_ (.I(_01013_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13599_ (.I(_01119_),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13600_ (.A1(_01120_),
    .A2(\register_file[11][0] ),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13601_ (.I(_01029_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13602_ (.I(_01122_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13603_ (.A1(_01123_),
    .A2(\register_file[10][0] ),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13604_ (.I(_01074_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13605_ (.I(_01125_),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13606_ (.A1(_01121_),
    .A2(_01124_),
    .B(_01126_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13607_ (.A1(_01118_),
    .A2(_01127_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13608_ (.I(_01017_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13609_ (.I(_01129_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13610_ (.A1(_01130_),
    .A2(\register_file[12][0] ),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13611_ (.I(_01034_),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13612_ (.I(_01132_),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13613_ (.I(_01037_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13614_ (.I(_01134_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13615_ (.A1(_01135_),
    .A2(\register_file[13][0] ),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13616_ (.A1(_01131_),
    .A2(_01133_),
    .A3(_01136_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13617_ (.I(_01029_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13618_ (.I(_01138_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13619_ (.A1(_01139_),
    .A2(\register_file[14][0] ),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13620_ (.I(_01093_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13621_ (.I(_01095_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13622_ (.I(_01142_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13623_ (.A1(_01143_),
    .A2(\register_file[15][0] ),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13624_ (.A1(_01140_),
    .A2(_01141_),
    .A3(_01144_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13625_ (.I(_01021_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13626_ (.I(_01146_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13627_ (.I(_01147_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13628_ (.A1(_01137_),
    .A2(_01145_),
    .A3(_01148_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13629_ (.A1(_01128_),
    .A2(_01149_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13630_ (.I(_01014_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13631_ (.I(_01151_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13632_ (.A1(_01152_),
    .A2(\register_file[6][0] ),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13633_ (.I(\register_file[7][0] ),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13634_ (.I(_01095_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13635_ (.I(_01155_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13636_ (.A1(_01154_),
    .A2(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13637_ (.I(_01023_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13638_ (.I(_01158_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13639_ (.A1(_01153_),
    .A2(_01157_),
    .A3(_01159_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13640_ (.I(_00993_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13641_ (.I(_01161_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13642_ (.I(\register_file[4][0] ),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13643_ (.A1(_01162_),
    .A2(_01163_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13644_ (.I(\register_file[5][0] ),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13645_ (.I(_00998_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13646_ (.I(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13647_ (.A1(_01165_),
    .A2(_01167_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13648_ (.I(_01033_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13649_ (.I(_01169_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13650_ (.A1(_01164_),
    .A2(_01168_),
    .A3(_01170_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13651_ (.A1(_01160_),
    .A2(_01171_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13652_ (.I(_01051_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13653_ (.A1(_01172_),
    .A2(_01173_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13654_ (.I(_01024_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13655_ (.I(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13656_ (.I(_01176_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _13657_ (.I(_00999_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _13658_ (.I(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13659_ (.A1(\register_file[2][0] ),
    .A2(_01179_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13660_ (.I(\register_file[3][0] ),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13661_ (.I(_01179_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13662_ (.A1(_01181_),
    .A2(_01182_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13663_ (.A1(_01177_),
    .A2(_01180_),
    .A3(_01183_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13664_ (.I(_01003_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13665_ (.I(_01185_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13666_ (.I(net9),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13667_ (.I(_01187_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13668_ (.A1(_01186_),
    .A2(\register_file[1][0] ),
    .B(_01188_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13669_ (.A1(_01184_),
    .A2(_01189_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13670_ (.I(_01190_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13671_ (.A1(_01174_),
    .A2(_01191_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13672_ (.I(net10),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13673_ (.I(_01193_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13674_ (.I(_01194_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13675_ (.A1(_01150_),
    .A2(_01192_),
    .A3(_01195_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13676_ (.A1(_01005_),
    .A2(_01030_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13677_ (.I(_01187_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _13678_ (.A1(_01197_),
    .A2(_01104_),
    .A3(_01198_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13679_ (.I(_01199_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13680_ (.I(_01200_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13681_ (.A1(_01106_),
    .A2(_01196_),
    .B(_01201_),
    .ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13682_ (.I(_00994_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13683_ (.A1(_01202_),
    .A2(\register_file[16][1] ),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13684_ (.A1(_01000_),
    .A2(\register_file[17][1] ),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13685_ (.A1(_01203_),
    .A2(_01204_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13686_ (.A1(_01205_),
    .A2(_01006_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13687_ (.A1(_01206_),
    .A2(_01011_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13688_ (.A1(_01015_),
    .A2(\register_file[19][1] ),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13689_ (.A1(_01019_),
    .A2(\register_file[18][1] ),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13690_ (.A1(_01208_),
    .A2(_01209_),
    .B(_01026_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13691_ (.A1(_01207_),
    .A2(_01210_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13692_ (.A1(_01031_),
    .A2(\register_file[20][1] ),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13693_ (.A1(_01039_),
    .A2(\register_file[21][1] ),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13694_ (.A1(_01212_),
    .A2(_01036_),
    .A3(_01213_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13695_ (.A1(_01043_),
    .A2(\register_file[22][1] ),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13696_ (.I(_01047_),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13697_ (.A1(_01216_),
    .A2(\register_file[23][1] ),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13698_ (.A1(_01215_),
    .A2(_01046_),
    .A3(_01217_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13699_ (.A1(_01214_),
    .A2(_01218_),
    .A3(_01052_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13700_ (.A1(_01211_),
    .A2(_01219_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13701_ (.A1(_01056_),
    .A2(\register_file[24][1] ),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13702_ (.A1(_01059_),
    .A2(\register_file[25][1] ),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13703_ (.A1(_01221_),
    .A2(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13704_ (.A1(_01223_),
    .A2(_01063_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13705_ (.I(_01065_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13706_ (.A1(_01224_),
    .A2(_01225_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13707_ (.A1(_01069_),
    .A2(\register_file[27][1] ),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13708_ (.A1(_01072_),
    .A2(\register_file[26][1] ),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13709_ (.A1(_01227_),
    .A2(_01228_),
    .B(_01076_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13710_ (.A1(_01226_),
    .A2(_01229_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13711_ (.A1(_01081_),
    .A2(\register_file[28][1] ),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13712_ (.A1(_01086_),
    .A2(\register_file[29][1] ),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13713_ (.A1(_01231_),
    .A2(_01084_),
    .A3(_01232_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13714_ (.A1(_01090_),
    .A2(\register_file[30][1] ),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13715_ (.A1(_01097_),
    .A2(\register_file[31][1] ),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13716_ (.A1(_01234_),
    .A2(_01094_),
    .A3(_01235_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13717_ (.I(_01100_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13718_ (.A1(_01233_),
    .A2(_01236_),
    .A3(_01237_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13719_ (.A1(_01230_),
    .A2(_01238_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13720_ (.A1(_01220_),
    .A2(_01239_),
    .A3(_01105_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13721_ (.A1(_01108_),
    .A2(\register_file[8][1] ),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13722_ (.I(_01110_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13723_ (.A1(_01242_),
    .A2(\register_file[9][1] ),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13724_ (.A1(_01241_),
    .A2(_01243_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13725_ (.A1(_01244_),
    .A2(_01115_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13726_ (.A1(_01245_),
    .A2(_01117_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13727_ (.I(_01119_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13728_ (.A1(_01247_),
    .A2(\register_file[11][1] ),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13729_ (.I(_01122_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13730_ (.A1(_01249_),
    .A2(\register_file[10][1] ),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13731_ (.A1(_01248_),
    .A2(_01250_),
    .B(_01126_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13732_ (.A1(_01246_),
    .A2(_01251_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13733_ (.I(_01129_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13734_ (.A1(_01253_),
    .A2(\register_file[12][1] ),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13735_ (.A1(_01135_),
    .A2(\register_file[13][1] ),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13736_ (.A1(_01254_),
    .A2(_01133_),
    .A3(_01255_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13737_ (.A1(_01139_),
    .A2(\register_file[14][1] ),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13738_ (.I(_01093_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13739_ (.A1(_01143_),
    .A2(\register_file[15][1] ),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13740_ (.A1(_01257_),
    .A2(_01258_),
    .A3(_01259_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13741_ (.A1(_01256_),
    .A2(_01260_),
    .A3(_01148_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13742_ (.A1(_01252_),
    .A2(_01261_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13743_ (.A1(_01152_),
    .A2(\register_file[6][1] ),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13744_ (.I(\register_file[7][1] ),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13745_ (.A1(_01264_),
    .A2(_01156_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13746_ (.I(_01158_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13747_ (.A1(_01263_),
    .A2(_01265_),
    .A3(_01266_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13748_ (.I(\register_file[4][1] ),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13749_ (.A1(_01162_),
    .A2(_01268_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13750_ (.I(\register_file[5][1] ),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13751_ (.I(_01166_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13752_ (.A1(_01270_),
    .A2(_01271_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13753_ (.I(_01169_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13754_ (.A1(_01269_),
    .A2(_01272_),
    .A3(_01273_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13755_ (.A1(_01267_),
    .A2(_01274_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13756_ (.A1(_01275_),
    .A2(_01173_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _13757_ (.I(_01178_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13758_ (.I(_01277_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13759_ (.A1(_01278_),
    .A2(\register_file[2][1] ),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13760_ (.I(\register_file[3][1] ),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13761_ (.A1(_01280_),
    .A2(_01182_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13762_ (.A1(_01177_),
    .A2(_01279_),
    .A3(_01281_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13763_ (.A1(_01186_),
    .A2(\register_file[1][1] ),
    .B(_01188_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13764_ (.A1(_01282_),
    .A2(_01283_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13765_ (.I(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13766_ (.A1(_01276_),
    .A2(_01285_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13767_ (.A1(_01262_),
    .A2(_01286_),
    .A3(_01195_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13768_ (.A1(_01240_),
    .A2(_01287_),
    .B(_01201_),
    .ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13769_ (.A1(_01202_),
    .A2(\register_file[16][2] ),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13770_ (.A1(_01000_),
    .A2(\register_file[17][2] ),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13771_ (.A1(_01288_),
    .A2(_01289_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13772_ (.A1(_01290_),
    .A2(_01006_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13773_ (.I(_01009_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13774_ (.A1(_01291_),
    .A2(_01292_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13775_ (.A1(_01015_),
    .A2(\register_file[19][2] ),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13776_ (.A1(_01019_),
    .A2(\register_file[18][2] ),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13777_ (.A1(_01294_),
    .A2(_01295_),
    .B(_01026_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13778_ (.A1(_01293_),
    .A2(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13779_ (.A1(_01031_),
    .A2(\register_file[20][2] ),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13780_ (.A1(_01039_),
    .A2(\register_file[21][2] ),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13781_ (.A1(_01298_),
    .A2(_01036_),
    .A3(_01299_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13782_ (.A1(_01043_),
    .A2(\register_file[22][2] ),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13783_ (.A1(_01216_),
    .A2(\register_file[23][2] ),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13784_ (.A1(_01301_),
    .A2(_01046_),
    .A3(_01302_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13785_ (.A1(_01300_),
    .A2(_01303_),
    .A3(_01052_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13786_ (.A1(_01297_),
    .A2(_01304_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13787_ (.A1(_01056_),
    .A2(\register_file[24][2] ),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13788_ (.I(_00998_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13789_ (.I(_01307_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13790_ (.A1(_01308_),
    .A2(\register_file[25][2] ),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13791_ (.A1(_01306_),
    .A2(_01309_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13792_ (.A1(_01310_),
    .A2(_01063_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13793_ (.A1(_01311_),
    .A2(_01225_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13794_ (.I(_01068_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13795_ (.A1(_01313_),
    .A2(\register_file[27][2] ),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13796_ (.A1(_01072_),
    .A2(\register_file[26][2] ),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13797_ (.A1(_01314_),
    .A2(_01315_),
    .B(_01076_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13798_ (.A1(_01312_),
    .A2(_01316_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13799_ (.I(_01017_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13800_ (.I(_01318_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13801_ (.A1(_01319_),
    .A2(\register_file[28][2] ),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13802_ (.A1(_01086_),
    .A2(\register_file[29][2] ),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13803_ (.A1(_01320_),
    .A2(_01084_),
    .A3(_01321_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13804_ (.I(_01089_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13805_ (.A1(_01323_),
    .A2(\register_file[30][2] ),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13806_ (.I(_01092_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13807_ (.I(_01325_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13808_ (.I(_01096_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13809_ (.A1(_01327_),
    .A2(\register_file[31][2] ),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13810_ (.A1(_01324_),
    .A2(_01326_),
    .A3(_01328_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13811_ (.A1(_01322_),
    .A2(_01329_),
    .A3(_01237_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13812_ (.A1(_01317_),
    .A2(_01330_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13813_ (.A1(_01305_),
    .A2(_01331_),
    .A3(_01105_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13814_ (.A1(_01108_),
    .A2(\register_file[8][2] ),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13815_ (.A1(_01242_),
    .A2(\register_file[9][2] ),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13816_ (.A1(_01333_),
    .A2(_01334_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13817_ (.A1(_01335_),
    .A2(_01115_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13818_ (.A1(_01336_),
    .A2(_01117_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13819_ (.A1(_01247_),
    .A2(\register_file[11][2] ),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13820_ (.A1(_01249_),
    .A2(\register_file[10][2] ),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13821_ (.A1(_01338_),
    .A2(_01339_),
    .B(_01126_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13822_ (.A1(_01337_),
    .A2(_01340_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13823_ (.A1(_01253_),
    .A2(\register_file[12][2] ),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13824_ (.I(_01132_),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13825_ (.I(_01134_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13826_ (.A1(_01344_),
    .A2(\register_file[13][2] ),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13827_ (.A1(_01342_),
    .A2(_01343_),
    .A3(_01345_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13828_ (.A1(_01139_),
    .A2(\register_file[14][2] ),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13829_ (.A1(_01143_),
    .A2(\register_file[15][2] ),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13830_ (.A1(_01347_),
    .A2(_01258_),
    .A3(_01348_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13831_ (.A1(_01346_),
    .A2(_01349_),
    .A3(_01148_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13832_ (.A1(_01341_),
    .A2(_01350_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13833_ (.A1(_01152_),
    .A2(\register_file[6][2] ),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13834_ (.I(\register_file[7][2] ),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13835_ (.I(_00998_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13836_ (.I(_01354_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13837_ (.A1(_01353_),
    .A2(_01355_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13838_ (.A1(_01352_),
    .A2(_01356_),
    .A3(_01266_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13839_ (.I(\register_file[4][2] ),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13840_ (.A1(_01162_),
    .A2(_01358_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13841_ (.I(\register_file[5][2] ),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13842_ (.A1(_01360_),
    .A2(_01271_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13843_ (.A1(_01359_),
    .A2(_01361_),
    .A3(_01273_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13844_ (.A1(_01357_),
    .A2(_01362_),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13845_ (.A1(_01363_),
    .A2(_01173_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13846_ (.A1(_01278_),
    .A2(\register_file[2][2] ),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13847_ (.I(\register_file[3][2] ),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13848_ (.A1(_01366_),
    .A2(_01182_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13849_ (.A1(_01177_),
    .A2(_01365_),
    .A3(_01367_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13850_ (.I(_01185_),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13851_ (.I(_01187_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13852_ (.I(_01370_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13853_ (.A1(_01369_),
    .A2(\register_file[1][2] ),
    .B(_01371_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13854_ (.A1(_01368_),
    .A2(_01372_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13855_ (.I(_01373_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13856_ (.A1(_01364_),
    .A2(_01374_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13857_ (.A1(_01351_),
    .A2(_01375_),
    .A3(_01195_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13858_ (.A1(_01332_),
    .A2(_01376_),
    .B(_01201_),
    .ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13859_ (.A1(_01202_),
    .A2(\register_file[16][3] ),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13860_ (.A1(_01000_),
    .A2(\register_file[17][3] ),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13861_ (.A1(_01377_),
    .A2(_01378_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13862_ (.A1(_01379_),
    .A2(_01006_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13863_ (.A1(_01380_),
    .A2(_01292_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13864_ (.I(_01014_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13865_ (.A1(_01382_),
    .A2(\register_file[19][3] ),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13866_ (.A1(_01019_),
    .A2(\register_file[18][3] ),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13867_ (.A1(_01383_),
    .A2(_01384_),
    .B(_01026_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13868_ (.A1(_01381_),
    .A2(_01385_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13869_ (.I(_01030_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13870_ (.A1(_01387_),
    .A2(\register_file[20][3] ),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13871_ (.A1(_01039_),
    .A2(\register_file[21][3] ),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13872_ (.A1(_01388_),
    .A2(_01036_),
    .A3(_01389_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13873_ (.A1(_01043_),
    .A2(\register_file[22][3] ),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13874_ (.A1(_01216_),
    .A2(\register_file[23][3] ),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13875_ (.A1(_01391_),
    .A2(_01046_),
    .A3(_01392_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13876_ (.I(_01146_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13877_ (.I(_01394_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13878_ (.A1(_01390_),
    .A2(_01393_),
    .A3(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13879_ (.A1(_01386_),
    .A2(_01396_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13880_ (.A1(_01056_),
    .A2(\register_file[24][3] ),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13881_ (.A1(_01308_),
    .A2(\register_file[25][3] ),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13882_ (.A1(_01398_),
    .A2(_01399_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13883_ (.A1(_01400_),
    .A2(_01063_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13884_ (.A1(_01401_),
    .A2(_01225_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13885_ (.A1(_01313_),
    .A2(\register_file[27][3] ),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13886_ (.I(_01029_),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13887_ (.I(_01404_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13888_ (.A1(_01405_),
    .A2(\register_file[26][3] ),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13889_ (.A1(_01403_),
    .A2(_01406_),
    .B(_01076_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13890_ (.A1(_01402_),
    .A2(_01407_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13891_ (.A1(_01319_),
    .A2(\register_file[28][3] ),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13892_ (.I(_01083_),
    .Z(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13893_ (.I(_01085_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13894_ (.A1(_01411_),
    .A2(\register_file[29][3] ),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13895_ (.A1(_01409_),
    .A2(_01410_),
    .A3(_01412_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13896_ (.A1(_01323_),
    .A2(\register_file[30][3] ),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13897_ (.A1(_01327_),
    .A2(\register_file[31][3] ),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13898_ (.A1(_01414_),
    .A2(_01326_),
    .A3(_01415_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13899_ (.A1(_01413_),
    .A2(_01416_),
    .A3(_01237_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13900_ (.A1(_01408_),
    .A2(_01417_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13901_ (.A1(_01397_),
    .A2(_01418_),
    .A3(_01105_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13902_ (.A1(_01108_),
    .A2(\register_file[8][3] ),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13903_ (.A1(_01242_),
    .A2(\register_file[9][3] ),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13904_ (.A1(_01420_),
    .A2(_01421_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13905_ (.I(_01004_),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13906_ (.I(_01423_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13907_ (.A1(_01422_),
    .A2(_01424_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13908_ (.I(net9),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13909_ (.I(_01426_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13910_ (.A1(_01425_),
    .A2(_01427_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13911_ (.A1(_01247_),
    .A2(\register_file[11][3] ),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13912_ (.A1(_01249_),
    .A2(\register_file[10][3] ),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13913_ (.I(_01125_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13914_ (.A1(_01429_),
    .A2(_01430_),
    .B(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13915_ (.A1(_01428_),
    .A2(_01432_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13916_ (.A1(_01253_),
    .A2(\register_file[12][3] ),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13917_ (.A1(_01344_),
    .A2(\register_file[13][3] ),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13918_ (.A1(_01434_),
    .A2(_01343_),
    .A3(_01435_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13919_ (.A1(_01139_),
    .A2(\register_file[14][3] ),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13920_ (.A1(_01143_),
    .A2(\register_file[15][3] ),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13921_ (.A1(_01437_),
    .A2(_01258_),
    .A3(_01438_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13922_ (.A1(_01436_),
    .A2(_01439_),
    .A3(_01148_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13923_ (.A1(_01433_),
    .A2(_01440_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13924_ (.A1(_01152_),
    .A2(\register_file[6][3] ),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13925_ (.I(\register_file[7][3] ),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13926_ (.A1(_01443_),
    .A2(_01355_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13927_ (.A1(_01442_),
    .A2(_01444_),
    .A3(_01266_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13928_ (.I(\register_file[4][3] ),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13929_ (.A1(_01162_),
    .A2(_01446_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13930_ (.I(\register_file[5][3] ),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13931_ (.A1(_01448_),
    .A2(_01271_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13932_ (.A1(_01447_),
    .A2(_01449_),
    .A3(_01273_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13933_ (.A1(_01445_),
    .A2(_01450_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13934_ (.A1(_01451_),
    .A2(_01173_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13935_ (.A1(_01278_),
    .A2(\register_file[2][3] ),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13936_ (.I(\register_file[3][3] ),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13937_ (.I(_01095_),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13938_ (.I(_01455_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13939_ (.A1(_01454_),
    .A2(_01456_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13940_ (.A1(_01177_),
    .A2(_01453_),
    .A3(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13941_ (.A1(_01369_),
    .A2(\register_file[1][3] ),
    .B(_01371_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13942_ (.A1(_01458_),
    .A2(_01459_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13943_ (.I(_01460_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13944_ (.A1(_01452_),
    .A2(_01461_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13945_ (.A1(_01441_),
    .A2(_01462_),
    .A3(_01195_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13946_ (.A1(_01419_),
    .A2(_01463_),
    .B(_01201_),
    .ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13947_ (.A1(_01202_),
    .A2(\register_file[24][4] ),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13948_ (.A1(_01000_),
    .A2(\register_file[25][4] ),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13949_ (.A1(_01464_),
    .A2(_01465_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13950_ (.A1(_01466_),
    .A2(_01006_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13951_ (.I(_01370_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13952_ (.A1(_01467_),
    .A2(_01468_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13953_ (.A1(_01382_),
    .A2(\register_file[27][4] ),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13954_ (.A1(_01019_),
    .A2(\register_file[26][4] ),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13955_ (.A1(_01470_),
    .A2(_01471_),
    .B(_01026_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13956_ (.A1(_01469_),
    .A2(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13957_ (.A1(_01387_),
    .A2(\register_file[28][4] ),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13958_ (.I(_01035_),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13959_ (.A1(_01039_),
    .A2(\register_file[29][4] ),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13960_ (.A1(_01474_),
    .A2(_01475_),
    .A3(_01476_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13961_ (.I(_01042_),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13962_ (.A1(_01478_),
    .A2(\register_file[30][4] ),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13963_ (.I(_01045_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13964_ (.A1(_01216_),
    .A2(\register_file[31][4] ),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13965_ (.A1(_01479_),
    .A2(_01480_),
    .A3(_01481_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13966_ (.A1(_01477_),
    .A2(_01482_),
    .A3(_01395_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13967_ (.A1(_01473_),
    .A2(_01483_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13968_ (.A1(_01056_),
    .A2(\register_file[16][4] ),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13969_ (.A1(_01308_),
    .A2(\register_file[17][4] ),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13970_ (.A1(_01485_),
    .A2(_01486_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13971_ (.I(_01062_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13972_ (.A1(_01487_),
    .A2(_01488_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13973_ (.I(_01009_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13974_ (.A1(_01489_),
    .A2(_01490_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13975_ (.A1(_01313_),
    .A2(\register_file[19][4] ),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13976_ (.A1(_01405_),
    .A2(\register_file[18][4] ),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13977_ (.I(_01075_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13978_ (.A1(_01492_),
    .A2(_01493_),
    .B(_01494_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13979_ (.A1(_01491_),
    .A2(_01495_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13980_ (.A1(_01319_),
    .A2(\register_file[20][4] ),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13981_ (.A1(_01411_),
    .A2(\register_file[21][4] ),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13982_ (.A1(_01497_),
    .A2(_01410_),
    .A3(_01498_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13983_ (.A1(_01323_),
    .A2(\register_file[22][4] ),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13984_ (.A1(_01327_),
    .A2(\register_file[23][4] ),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13985_ (.A1(_01500_),
    .A2(_01326_),
    .A3(_01501_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13986_ (.A1(_01499_),
    .A2(_01502_),
    .A3(_01237_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13987_ (.A1(_01496_),
    .A2(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13988_ (.I(net10),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13989_ (.I(_01505_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13990_ (.A1(_01484_),
    .A2(_01504_),
    .A3(_01506_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13991_ (.I(_01107_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13992_ (.A1(_01508_),
    .A2(\register_file[8][4] ),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13993_ (.A1(_01242_),
    .A2(\register_file[9][4] ),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13994_ (.A1(_01509_),
    .A2(_01510_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13995_ (.A1(_01511_),
    .A2(_01424_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13996_ (.A1(_01512_),
    .A2(_01427_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13997_ (.A1(_01247_),
    .A2(\register_file[11][4] ),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13998_ (.A1(_01249_),
    .A2(\register_file[10][4] ),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13999_ (.A1(_01514_),
    .A2(_01515_),
    .B(_01431_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14000_ (.A1(_01513_),
    .A2(_01516_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14001_ (.A1(_01253_),
    .A2(\register_file[12][4] ),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14002_ (.A1(_01344_),
    .A2(\register_file[13][4] ),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14003_ (.A1(_01518_),
    .A2(_01343_),
    .A3(_01519_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14004_ (.A1(_01139_),
    .A2(\register_file[14][4] ),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14005_ (.A1(_01143_),
    .A2(\register_file[15][4] ),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14006_ (.A1(_01521_),
    .A2(_01258_),
    .A3(_01522_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14007_ (.A1(_01520_),
    .A2(_01523_),
    .A3(_01148_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14008_ (.A1(_01517_),
    .A2(_01524_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14009_ (.A1(_01152_),
    .A2(\register_file[6][4] ),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14010_ (.I(\register_file[7][4] ),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14011_ (.A1(_01527_),
    .A2(_01355_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14012_ (.A1(_01526_),
    .A2(_01528_),
    .A3(_01266_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14013_ (.I(_00993_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14014_ (.I(_01530_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14015_ (.I(\register_file[4][4] ),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14016_ (.A1(_01531_),
    .A2(_01532_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14017_ (.I(\register_file[5][4] ),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14018_ (.A1(_01534_),
    .A2(_01271_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14019_ (.A1(_01533_),
    .A2(_01535_),
    .A3(_01273_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14020_ (.A1(_01529_),
    .A2(_01536_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14021_ (.I(_01146_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14022_ (.A1(_01537_),
    .A2(_01538_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14023_ (.A1(_01278_),
    .A2(\register_file[2][4] ),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14024_ (.I(\register_file[3][4] ),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14025_ (.A1(_01541_),
    .A2(_01456_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14026_ (.A1(_01177_),
    .A2(_01540_),
    .A3(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14027_ (.A1(_01369_),
    .A2(\register_file[1][4] ),
    .B(_01371_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14028_ (.A1(_01543_),
    .A2(_01544_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14029_ (.I(_01545_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14030_ (.A1(_01539_),
    .A2(_01546_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14031_ (.A1(_01525_),
    .A2(_01547_),
    .A3(_01195_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14032_ (.A1(_01507_),
    .A2(_01548_),
    .B(_01201_),
    .ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14033_ (.A1(_01202_),
    .A2(\register_file[24][5] ),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14034_ (.I(_00999_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14035_ (.A1(_01550_),
    .A2(\register_file[25][5] ),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14036_ (.A1(_01549_),
    .A2(_01551_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14037_ (.I(_01005_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14038_ (.A1(_01552_),
    .A2(_01553_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14039_ (.A1(_01554_),
    .A2(_01468_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14040_ (.A1(_01382_),
    .A2(\register_file[27][5] ),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14041_ (.I(_01018_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14042_ (.A1(_01557_),
    .A2(\register_file[26][5] ),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14043_ (.I(_01074_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14044_ (.I(_01559_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14045_ (.A1(_01556_),
    .A2(_01558_),
    .B(_01560_),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14046_ (.A1(_01555_),
    .A2(_01561_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14047_ (.A1(_01387_),
    .A2(\register_file[28][5] ),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14048_ (.I(_01038_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14049_ (.A1(_01564_),
    .A2(\register_file[29][5] ),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14050_ (.A1(_01563_),
    .A2(_01475_),
    .A3(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14051_ (.A1(_01478_),
    .A2(\register_file[30][5] ),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14052_ (.A1(_01216_),
    .A2(\register_file[31][5] ),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14053_ (.A1(_01567_),
    .A2(_01480_),
    .A3(_01568_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14054_ (.A1(_01566_),
    .A2(_01569_),
    .A3(_01395_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14055_ (.A1(_01562_),
    .A2(_01570_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14056_ (.I(_01055_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14057_ (.A1(_01572_),
    .A2(\register_file[16][5] ),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14058_ (.A1(_01308_),
    .A2(\register_file[17][5] ),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14059_ (.A1(_01573_),
    .A2(_01574_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14060_ (.A1(_01575_),
    .A2(_01488_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14061_ (.A1(_01576_),
    .A2(_01490_),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14062_ (.A1(_01313_),
    .A2(\register_file[19][5] ),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14063_ (.A1(_01405_),
    .A2(\register_file[18][5] ),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14064_ (.A1(_01578_),
    .A2(_01579_),
    .B(_01494_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14065_ (.A1(_01577_),
    .A2(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14066_ (.A1(_01319_),
    .A2(\register_file[20][5] ),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14067_ (.A1(_01411_),
    .A2(\register_file[21][5] ),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14068_ (.A1(_01582_),
    .A2(_01410_),
    .A3(_01583_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14069_ (.A1(_01323_),
    .A2(\register_file[22][5] ),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14070_ (.A1(_01327_),
    .A2(\register_file[23][5] ),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14071_ (.A1(_01585_),
    .A2(_01326_),
    .A3(_01586_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14072_ (.A1(_01584_),
    .A2(_01587_),
    .A3(_01237_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14073_ (.A1(_01581_),
    .A2(_01588_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14074_ (.A1(_01571_),
    .A2(_01589_),
    .A3(_01506_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14075_ (.A1(_01508_),
    .A2(\register_file[8][5] ),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14076_ (.A1(_01242_),
    .A2(\register_file[9][5] ),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14077_ (.A1(_01591_),
    .A2(_01592_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14078_ (.A1(_01593_),
    .A2(_01424_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14079_ (.A1(_01594_),
    .A2(_01427_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14080_ (.A1(_01247_),
    .A2(\register_file[11][5] ),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14081_ (.A1(_01249_),
    .A2(\register_file[10][5] ),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14082_ (.A1(_01596_),
    .A2(_01597_),
    .B(_01431_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14083_ (.A1(_01595_),
    .A2(_01598_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14084_ (.A1(_01253_),
    .A2(\register_file[12][5] ),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14085_ (.A1(_01344_),
    .A2(\register_file[13][5] ),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14086_ (.A1(_01600_),
    .A2(_01343_),
    .A3(_01601_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14087_ (.I(_01138_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14088_ (.A1(_01603_),
    .A2(\register_file[14][5] ),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14089_ (.I(_01142_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14090_ (.A1(_01605_),
    .A2(\register_file[15][5] ),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14091_ (.A1(_01604_),
    .A2(_01258_),
    .A3(_01606_),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14092_ (.I(_01147_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14093_ (.A1(_01602_),
    .A2(_01607_),
    .A3(_01608_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14094_ (.A1(_01599_),
    .A2(_01609_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14095_ (.I(_01151_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14096_ (.A1(_01611_),
    .A2(\register_file[6][5] ),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14097_ (.I(\register_file[7][5] ),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14098_ (.A1(_01613_),
    .A2(_01355_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14099_ (.A1(_01612_),
    .A2(_01614_),
    .A3(_01266_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14100_ (.I(\register_file[4][5] ),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14101_ (.A1(_01531_),
    .A2(_01616_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14102_ (.I(\register_file[5][5] ),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14103_ (.A1(_01618_),
    .A2(_01271_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14104_ (.A1(_01617_),
    .A2(_01619_),
    .A3(_01273_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14105_ (.A1(_01615_),
    .A2(_01620_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14106_ (.A1(_01621_),
    .A2(_01538_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14107_ (.I(_01176_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14108_ (.A1(_01278_),
    .A2(\register_file[2][5] ),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14109_ (.I(\register_file[3][5] ),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14110_ (.A1(_01625_),
    .A2(_01456_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14111_ (.A1(_01623_),
    .A2(_01624_),
    .A3(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14112_ (.A1(_01369_),
    .A2(\register_file[1][5] ),
    .B(_01371_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14113_ (.A1(_01627_),
    .A2(_01628_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14114_ (.I(_01629_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14115_ (.A1(_01622_),
    .A2(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14116_ (.I(_01194_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14117_ (.A1(_01610_),
    .A2(_01631_),
    .A3(_01632_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14118_ (.I(_01200_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14119_ (.A1(_01590_),
    .A2(_01633_),
    .B(_01634_),
    .ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14120_ (.I(_00994_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14121_ (.A1(_01635_),
    .A2(\register_file[24][6] ),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14122_ (.A1(_01550_),
    .A2(\register_file[25][6] ),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14123_ (.A1(_01636_),
    .A2(_01637_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14124_ (.A1(_01638_),
    .A2(_01553_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14125_ (.A1(_01639_),
    .A2(_01468_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14126_ (.A1(_01382_),
    .A2(\register_file[27][6] ),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14127_ (.A1(_01557_),
    .A2(\register_file[26][6] ),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14128_ (.A1(_01641_),
    .A2(_01642_),
    .B(_01560_),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14129_ (.A1(_01640_),
    .A2(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14130_ (.A1(_01387_),
    .A2(\register_file[28][6] ),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14131_ (.A1(_01564_),
    .A2(\register_file[29][6] ),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14132_ (.A1(_01645_),
    .A2(_01475_),
    .A3(_01646_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14133_ (.A1(_01478_),
    .A2(\register_file[30][6] ),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14134_ (.I(_01095_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14135_ (.I(_01649_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14136_ (.A1(_01650_),
    .A2(\register_file[31][6] ),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14137_ (.A1(_01648_),
    .A2(_01480_),
    .A3(_01651_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14138_ (.A1(_01647_),
    .A2(_01652_),
    .A3(_01395_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14139_ (.A1(_01644_),
    .A2(_01653_),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14140_ (.A1(_01572_),
    .A2(\register_file[16][6] ),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14141_ (.A1(_01308_),
    .A2(\register_file[17][6] ),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14142_ (.A1(_01655_),
    .A2(_01656_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14143_ (.A1(_01657_),
    .A2(_01488_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14144_ (.A1(_01658_),
    .A2(_01490_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14145_ (.A1(_01313_),
    .A2(\register_file[19][6] ),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14146_ (.A1(_01405_),
    .A2(\register_file[18][6] ),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14147_ (.A1(_01660_),
    .A2(_01661_),
    .B(_01494_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14148_ (.A1(_01659_),
    .A2(_01662_),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14149_ (.A1(_01319_),
    .A2(\register_file[20][6] ),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14150_ (.A1(_01411_),
    .A2(\register_file[21][6] ),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14151_ (.A1(_01664_),
    .A2(_01410_),
    .A3(_01665_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14152_ (.A1(_01323_),
    .A2(\register_file[22][6] ),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14153_ (.A1(_01327_),
    .A2(\register_file[23][6] ),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14154_ (.A1(_01667_),
    .A2(_01326_),
    .A3(_01668_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14155_ (.I(_01051_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14156_ (.I(_01670_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14157_ (.A1(_01666_),
    .A2(_01669_),
    .A3(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14158_ (.A1(_01663_),
    .A2(_01672_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14159_ (.A1(_01654_),
    .A2(_01673_),
    .A3(_01506_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14160_ (.A1(_01508_),
    .A2(\register_file[8][6] ),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14161_ (.I(_01110_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14162_ (.A1(_01676_),
    .A2(\register_file[9][6] ),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14163_ (.A1(_01675_),
    .A2(_01677_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14164_ (.A1(_01678_),
    .A2(_01424_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14165_ (.A1(_01679_),
    .A2(_01427_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14166_ (.I(_01037_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14167_ (.I(_01681_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14168_ (.A1(_01682_),
    .A2(\register_file[11][6] ),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14169_ (.I(_01122_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14170_ (.A1(_01684_),
    .A2(\register_file[10][6] ),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14171_ (.A1(_01683_),
    .A2(_01685_),
    .B(_01431_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14172_ (.A1(_01680_),
    .A2(_01686_),
    .ZN(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14173_ (.I(_01129_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14174_ (.A1(_01688_),
    .A2(\register_file[12][6] ),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14175_ (.A1(_01344_),
    .A2(\register_file[13][6] ),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14176_ (.A1(_01689_),
    .A2(_01343_),
    .A3(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14177_ (.A1(_01603_),
    .A2(\register_file[14][6] ),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14178_ (.I(_01092_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14179_ (.I(_01693_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14180_ (.A1(_01605_),
    .A2(\register_file[15][6] ),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14181_ (.A1(_01692_),
    .A2(_01694_),
    .A3(_01695_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14182_ (.A1(_01691_),
    .A2(_01696_),
    .A3(_01608_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14183_ (.A1(_01687_),
    .A2(_01697_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14184_ (.A1(_01611_),
    .A2(\register_file[6][6] ),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14185_ (.I(\register_file[7][6] ),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14186_ (.A1(_01700_),
    .A2(_01355_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14187_ (.I(_01158_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14188_ (.A1(_01699_),
    .A2(_01701_),
    .A3(_01702_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14189_ (.I(\register_file[4][6] ),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14190_ (.A1(_01531_),
    .A2(_01704_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14191_ (.I(\register_file[5][6] ),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14192_ (.I(_01166_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14193_ (.A1(_01706_),
    .A2(_01707_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14194_ (.I(_01169_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14195_ (.A1(_01705_),
    .A2(_01708_),
    .A3(_01709_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14196_ (.A1(_01703_),
    .A2(_01710_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14197_ (.A1(_01711_),
    .A2(_01538_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _14198_ (.I(_01277_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14199_ (.A1(_01713_),
    .A2(\register_file[2][6] ),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14200_ (.I(\register_file[3][6] ),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14201_ (.A1(_01715_),
    .A2(_01456_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14202_ (.A1(_01623_),
    .A2(_01714_),
    .A3(_01716_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14203_ (.A1(_01369_),
    .A2(\register_file[1][6] ),
    .B(_01371_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14204_ (.A1(_01717_),
    .A2(_01718_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14205_ (.I(_01719_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14206_ (.A1(_01712_),
    .A2(_01720_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14207_ (.A1(_01698_),
    .A2(_01721_),
    .A3(_01632_),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14208_ (.A1(_01674_),
    .A2(_01722_),
    .B(_01634_),
    .ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14209_ (.A1(_01635_),
    .A2(\register_file[24][7] ),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14210_ (.A1(_01550_),
    .A2(\register_file[25][7] ),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14211_ (.A1(_01723_),
    .A2(_01724_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14212_ (.A1(_01725_),
    .A2(_01553_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14213_ (.A1(_01726_),
    .A2(_01468_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14214_ (.A1(_01382_),
    .A2(\register_file[27][7] ),
    .ZN(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14215_ (.A1(_01557_),
    .A2(\register_file[26][7] ),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14216_ (.A1(_01728_),
    .A2(_01729_),
    .B(_01560_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14217_ (.A1(_01727_),
    .A2(_01730_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14218_ (.A1(_01387_),
    .A2(\register_file[28][7] ),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14219_ (.A1(_01564_),
    .A2(\register_file[29][7] ),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14220_ (.A1(_01732_),
    .A2(_01475_),
    .A3(_01733_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14221_ (.A1(_01478_),
    .A2(\register_file[30][7] ),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14222_ (.A1(_01650_),
    .A2(\register_file[31][7] ),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14223_ (.A1(_01735_),
    .A2(_01480_),
    .A3(_01736_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14224_ (.A1(_01734_),
    .A2(_01737_),
    .A3(_01395_),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14225_ (.A1(_01731_),
    .A2(_01738_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14226_ (.A1(_01572_),
    .A2(\register_file[16][7] ),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14227_ (.I(_01307_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14228_ (.A1(_01741_),
    .A2(\register_file[17][7] ),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14229_ (.A1(_01740_),
    .A2(_01742_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14230_ (.A1(_01743_),
    .A2(_01488_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14231_ (.A1(_01744_),
    .A2(_01490_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14232_ (.I(_01068_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14233_ (.A1(_01746_),
    .A2(\register_file[19][7] ),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14234_ (.A1(_01405_),
    .A2(\register_file[18][7] ),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14235_ (.A1(_01747_),
    .A2(_01748_),
    .B(_01494_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14236_ (.A1(_01745_),
    .A2(_01749_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14237_ (.I(_01318_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14238_ (.A1(_01751_),
    .A2(\register_file[20][7] ),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14239_ (.A1(_01411_),
    .A2(\register_file[21][7] ),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14240_ (.A1(_01752_),
    .A2(_01410_),
    .A3(_01753_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14241_ (.I(_01089_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14242_ (.A1(_01755_),
    .A2(\register_file[22][7] ),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14243_ (.I(_01325_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14244_ (.I(_01096_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14245_ (.A1(_01758_),
    .A2(\register_file[23][7] ),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14246_ (.A1(_01756_),
    .A2(_01757_),
    .A3(_01759_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14247_ (.A1(_01754_),
    .A2(_01760_),
    .A3(_01671_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14248_ (.A1(_01750_),
    .A2(_01761_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14249_ (.A1(_01739_),
    .A2(_01762_),
    .A3(_01506_),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14250_ (.A1(_01508_),
    .A2(\register_file[8][7] ),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14251_ (.A1(_01676_),
    .A2(\register_file[9][7] ),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14252_ (.A1(_01764_),
    .A2(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14253_ (.A1(_01766_),
    .A2(_01424_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14254_ (.A1(_01767_),
    .A2(_01427_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14255_ (.A1(_01682_),
    .A2(\register_file[11][7] ),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14256_ (.A1(_01684_),
    .A2(\register_file[10][7] ),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14257_ (.A1(_01769_),
    .A2(_01770_),
    .B(_01431_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14258_ (.A1(_01768_),
    .A2(_01771_),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14259_ (.A1(_01688_),
    .A2(\register_file[12][7] ),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14260_ (.I(_01033_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14261_ (.I(_01774_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14262_ (.I(_01134_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14263_ (.A1(_01776_),
    .A2(\register_file[13][7] ),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14264_ (.A1(_01773_),
    .A2(_01775_),
    .A3(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14265_ (.A1(_01603_),
    .A2(\register_file[14][7] ),
    .ZN(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14266_ (.A1(_01605_),
    .A2(\register_file[15][7] ),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14267_ (.A1(_01779_),
    .A2(_01694_),
    .A3(_01780_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14268_ (.A1(_01778_),
    .A2(_01781_),
    .A3(_01608_),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14269_ (.A1(_01772_),
    .A2(_01782_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14270_ (.A1(_01611_),
    .A2(\register_file[6][7] ),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14271_ (.I(\register_file[7][7] ),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14272_ (.I(_01354_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14273_ (.A1(_01785_),
    .A2(_01786_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14274_ (.A1(_01784_),
    .A2(_01787_),
    .A3(_01702_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14275_ (.I(\register_file[4][7] ),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14276_ (.A1(_01531_),
    .A2(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14277_ (.I(\register_file[5][7] ),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14278_ (.A1(_01791_),
    .A2(_01707_),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14279_ (.A1(_01790_),
    .A2(_01792_),
    .A3(_01709_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14280_ (.A1(_01788_),
    .A2(_01793_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14281_ (.A1(_01794_),
    .A2(_01538_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14282_ (.A1(_01713_),
    .A2(\register_file[2][7] ),
    .Z(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14283_ (.I(\register_file[3][7] ),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14284_ (.A1(_01797_),
    .A2(_01456_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14285_ (.A1(_01623_),
    .A2(_01796_),
    .A3(_01798_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14286_ (.I(_01185_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14287_ (.I(_01370_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14288_ (.A1(_01800_),
    .A2(\register_file[1][7] ),
    .B(_01801_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14289_ (.A1(_01799_),
    .A2(_01802_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14290_ (.I(_01803_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14291_ (.A1(_01795_),
    .A2(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14292_ (.A1(_01783_),
    .A2(_01805_),
    .A3(_01632_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14293_ (.A1(_01763_),
    .A2(_01806_),
    .B(_01634_),
    .ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14294_ (.A1(_01635_),
    .A2(\register_file[24][8] ),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14295_ (.A1(_01550_),
    .A2(\register_file[25][8] ),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14296_ (.A1(_01807_),
    .A2(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14297_ (.A1(_01809_),
    .A2(_01553_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14298_ (.I(_01187_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14299_ (.A1(_01810_),
    .A2(_01811_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14300_ (.I(_01014_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14301_ (.A1(_01813_),
    .A2(\register_file[27][8] ),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14302_ (.A1(_01557_),
    .A2(\register_file[26][8] ),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14303_ (.A1(_01814_),
    .A2(_01815_),
    .B(_01560_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14304_ (.A1(_01812_),
    .A2(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14305_ (.I(_01080_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14306_ (.A1(_01818_),
    .A2(\register_file[28][8] ),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14307_ (.A1(_01564_),
    .A2(\register_file[29][8] ),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14308_ (.A1(_01819_),
    .A2(_01475_),
    .A3(_01820_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14309_ (.A1(_01478_),
    .A2(\register_file[30][8] ),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14310_ (.A1(_01650_),
    .A2(\register_file[31][8] ),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14311_ (.A1(_01822_),
    .A2(_01480_),
    .A3(_01823_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14312_ (.I(_01394_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14313_ (.A1(_01821_),
    .A2(_01824_),
    .A3(_01825_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14314_ (.A1(_01817_),
    .A2(_01826_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14315_ (.A1(_01572_),
    .A2(\register_file[16][8] ),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14316_ (.A1(_01741_),
    .A2(\register_file[17][8] ),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14317_ (.A1(_01828_),
    .A2(_01829_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14318_ (.A1(_01830_),
    .A2(_01488_),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14319_ (.I(_01009_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14320_ (.A1(_01831_),
    .A2(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14321_ (.A1(_01746_),
    .A2(\register_file[19][8] ),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14322_ (.I(_01404_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14323_ (.A1(_01835_),
    .A2(\register_file[18][8] ),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14324_ (.A1(_01834_),
    .A2(_01836_),
    .B(_01494_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14325_ (.A1(_01833_),
    .A2(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14326_ (.A1(_01751_),
    .A2(\register_file[20][8] ),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14327_ (.I(_01083_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14328_ (.I(_01085_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14329_ (.A1(_01841_),
    .A2(\register_file[21][8] ),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14330_ (.A1(_01839_),
    .A2(_01840_),
    .A3(_01842_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14331_ (.A1(_01755_),
    .A2(\register_file[22][8] ),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14332_ (.A1(_01758_),
    .A2(\register_file[23][8] ),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14333_ (.A1(_01844_),
    .A2(_01757_),
    .A3(_01845_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14334_ (.A1(_01843_),
    .A2(_01846_),
    .A3(_01671_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14335_ (.A1(_01838_),
    .A2(_01847_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14336_ (.A1(_01827_),
    .A2(_01848_),
    .A3(_01506_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14337_ (.A1(_01508_),
    .A2(\register_file[8][8] ),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14338_ (.A1(_01676_),
    .A2(\register_file[9][8] ),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14339_ (.A1(_01850_),
    .A2(_01851_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14340_ (.I(_01423_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14341_ (.A1(_01852_),
    .A2(_01853_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14342_ (.I(_01426_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14343_ (.A1(_01854_),
    .A2(_01855_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14344_ (.A1(_01682_),
    .A2(\register_file[11][8] ),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14345_ (.A1(_01684_),
    .A2(\register_file[10][8] ),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14346_ (.I(_01125_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14347_ (.A1(_01857_),
    .A2(_01858_),
    .B(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14348_ (.A1(_01856_),
    .A2(_01860_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14349_ (.A1(_01688_),
    .A2(\register_file[12][8] ),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14350_ (.A1(_01776_),
    .A2(\register_file[13][8] ),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14351_ (.A1(_01862_),
    .A2(_01775_),
    .A3(_01863_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14352_ (.A1(_01603_),
    .A2(\register_file[14][8] ),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14353_ (.A1(_01605_),
    .A2(\register_file[15][8] ),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14354_ (.A1(_01865_),
    .A2(_01694_),
    .A3(_01866_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14355_ (.A1(_01864_),
    .A2(_01867_),
    .A3(_01608_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14356_ (.A1(_01861_),
    .A2(_01868_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14357_ (.A1(_01611_),
    .A2(\register_file[6][8] ),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14358_ (.I(\register_file[7][8] ),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14359_ (.A1(_01871_),
    .A2(_01786_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14360_ (.A1(_01870_),
    .A2(_01872_),
    .A3(_01702_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14361_ (.I(\register_file[4][8] ),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14362_ (.A1(_01531_),
    .A2(_01874_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14363_ (.I(\register_file[5][8] ),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14364_ (.A1(_01876_),
    .A2(_01707_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14365_ (.A1(_01875_),
    .A2(_01877_),
    .A3(_01709_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14366_ (.A1(_01873_),
    .A2(_01878_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14367_ (.A1(_01879_),
    .A2(_01538_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14368_ (.A1(_01713_),
    .A2(\register_file[2][8] ),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14369_ (.I(\register_file[3][8] ),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14370_ (.I(_01155_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14371_ (.A1(_01882_),
    .A2(_01883_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14372_ (.A1(_01623_),
    .A2(_01881_),
    .A3(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14373_ (.A1(_01800_),
    .A2(\register_file[1][8] ),
    .B(_01801_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14374_ (.A1(_01885_),
    .A2(_01886_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14375_ (.I(_01887_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14376_ (.A1(_01880_),
    .A2(_01888_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14377_ (.A1(_01869_),
    .A2(_01889_),
    .A3(_01632_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14378_ (.A1(_01849_),
    .A2(_01890_),
    .B(_01634_),
    .ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14379_ (.A1(_01635_),
    .A2(\register_file[24][9] ),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14380_ (.A1(_01550_),
    .A2(\register_file[25][9] ),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14381_ (.A1(_01891_),
    .A2(_01892_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14382_ (.A1(_01893_),
    .A2(_01553_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14383_ (.A1(_01894_),
    .A2(_01811_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14384_ (.A1(_01813_),
    .A2(\register_file[27][9] ),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14385_ (.A1(_01557_),
    .A2(\register_file[26][9] ),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14386_ (.A1(_01896_),
    .A2(_01897_),
    .B(_01560_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14387_ (.A1(_01895_),
    .A2(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14388_ (.A1(_01818_),
    .A2(\register_file[28][9] ),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14389_ (.I(_01035_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14390_ (.A1(_01564_),
    .A2(\register_file[29][9] ),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14391_ (.A1(_01900_),
    .A2(_01901_),
    .A3(_01902_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14392_ (.I(_01071_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14393_ (.A1(_01904_),
    .A2(\register_file[30][9] ),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14394_ (.I(_01045_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14395_ (.A1(_01650_),
    .A2(\register_file[31][9] ),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14396_ (.A1(_01905_),
    .A2(_01906_),
    .A3(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14397_ (.A1(_01903_),
    .A2(_01908_),
    .A3(_01825_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14398_ (.A1(_01899_),
    .A2(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14399_ (.A1(_01572_),
    .A2(\register_file[16][9] ),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14400_ (.A1(_01741_),
    .A2(\register_file[17][9] ),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14401_ (.A1(_01911_),
    .A2(_01912_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14402_ (.I(_01114_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14403_ (.A1(_01913_),
    .A2(_01914_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14404_ (.A1(_01915_),
    .A2(_01832_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14405_ (.A1(_01746_),
    .A2(\register_file[19][9] ),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14406_ (.A1(_01835_),
    .A2(\register_file[18][9] ),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14407_ (.I(_01075_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14408_ (.A1(_01917_),
    .A2(_01918_),
    .B(_01919_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14409_ (.A1(_01916_),
    .A2(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14410_ (.A1(_01751_),
    .A2(\register_file[20][9] ),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14411_ (.A1(_01841_),
    .A2(\register_file[21][9] ),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14412_ (.A1(_01922_),
    .A2(_01840_),
    .A3(_01923_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14413_ (.A1(_01755_),
    .A2(\register_file[22][9] ),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14414_ (.A1(_01758_),
    .A2(\register_file[23][9] ),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14415_ (.A1(_01925_),
    .A2(_01757_),
    .A3(_01926_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14416_ (.A1(_01924_),
    .A2(_01927_),
    .A3(_01671_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14417_ (.A1(_01921_),
    .A2(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14418_ (.I(_01505_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14419_ (.A1(_01910_),
    .A2(_01929_),
    .A3(_01930_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14420_ (.I(_01079_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14421_ (.A1(_01932_),
    .A2(\register_file[8][9] ),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14422_ (.A1(_01676_),
    .A2(\register_file[9][9] ),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14423_ (.A1(_01933_),
    .A2(_01934_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14424_ (.A1(_01935_),
    .A2(_01853_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14425_ (.A1(_01936_),
    .A2(_01855_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14426_ (.A1(_01682_),
    .A2(\register_file[11][9] ),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14427_ (.A1(_01684_),
    .A2(\register_file[10][9] ),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14428_ (.A1(_01938_),
    .A2(_01939_),
    .B(_01859_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14429_ (.A1(_01937_),
    .A2(_01940_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14430_ (.A1(_01688_),
    .A2(\register_file[12][9] ),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14431_ (.A1(_01776_),
    .A2(\register_file[13][9] ),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14432_ (.A1(_01942_),
    .A2(_01775_),
    .A3(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14433_ (.A1(_01603_),
    .A2(\register_file[14][9] ),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14434_ (.A1(_01605_),
    .A2(\register_file[15][9] ),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14435_ (.A1(_01945_),
    .A2(_01694_),
    .A3(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14436_ (.A1(_01944_),
    .A2(_01947_),
    .A3(_01608_),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14437_ (.A1(_01941_),
    .A2(_01948_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14438_ (.A1(_01611_),
    .A2(\register_file[6][9] ),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14439_ (.I(\register_file[7][9] ),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14440_ (.A1(_01951_),
    .A2(_01786_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14441_ (.A1(_01950_),
    .A2(_01952_),
    .A3(_01702_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14442_ (.I(_01530_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14443_ (.I(\register_file[4][9] ),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14444_ (.A1(_01954_),
    .A2(_01955_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14445_ (.I(\register_file[5][9] ),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14446_ (.A1(_01957_),
    .A2(_01707_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14447_ (.A1(_01956_),
    .A2(_01958_),
    .A3(_01709_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14448_ (.A1(_01953_),
    .A2(_01959_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14449_ (.I(_01146_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14450_ (.A1(_01960_),
    .A2(_01961_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14451_ (.A1(_01713_),
    .A2(\register_file[2][9] ),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14452_ (.I(\register_file[3][9] ),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14453_ (.A1(_01964_),
    .A2(_01883_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14454_ (.A1(_01623_),
    .A2(_01963_),
    .A3(_01965_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14455_ (.A1(_01800_),
    .A2(\register_file[1][9] ),
    .B(_01801_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14456_ (.A1(_01966_),
    .A2(_01967_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14457_ (.I(_01968_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14458_ (.A1(_01962_),
    .A2(_01969_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14459_ (.A1(_01949_),
    .A2(_01970_),
    .A3(_01632_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14460_ (.A1(_01931_),
    .A2(_01971_),
    .B(_01634_),
    .ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14461_ (.A1(_01635_),
    .A2(\register_file[24][10] ),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14462_ (.I(_01058_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14463_ (.A1(_01973_),
    .A2(\register_file[25][10] ),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14464_ (.A1(_01972_),
    .A2(_01974_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14465_ (.I(_01005_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14466_ (.A1(_01975_),
    .A2(_01976_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14467_ (.A1(_01977_),
    .A2(_01811_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14468_ (.A1(_01813_),
    .A2(\register_file[27][10] ),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14469_ (.I(_01018_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14470_ (.A1(_01980_),
    .A2(\register_file[26][10] ),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14471_ (.I(_01559_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14472_ (.A1(_01979_),
    .A2(_01981_),
    .B(_01982_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14473_ (.A1(_01978_),
    .A2(_01983_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14474_ (.A1(_01818_),
    .A2(\register_file[28][10] ),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14475_ (.I(_01038_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14476_ (.A1(_01986_),
    .A2(\register_file[29][10] ),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14477_ (.A1(_01985_),
    .A2(_01901_),
    .A3(_01987_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14478_ (.A1(_01904_),
    .A2(\register_file[30][10] ),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14479_ (.A1(_01650_),
    .A2(\register_file[31][10] ),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14480_ (.A1(_01989_),
    .A2(_01906_),
    .A3(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14481_ (.A1(_01988_),
    .A2(_01991_),
    .A3(_01825_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14482_ (.A1(_01984_),
    .A2(_01992_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14483_ (.I(_01055_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14484_ (.A1(_01994_),
    .A2(\register_file[16][10] ),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14485_ (.A1(_01741_),
    .A2(\register_file[17][10] ),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14486_ (.A1(_01995_),
    .A2(_01996_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14487_ (.A1(_01997_),
    .A2(_01914_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14488_ (.A1(_01998_),
    .A2(_01832_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14489_ (.A1(_01746_),
    .A2(\register_file[19][10] ),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14490_ (.A1(_01835_),
    .A2(\register_file[18][10] ),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14491_ (.A1(_02000_),
    .A2(_02001_),
    .B(_01919_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14492_ (.A1(_01999_),
    .A2(_02002_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14493_ (.A1(_01751_),
    .A2(\register_file[20][10] ),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14494_ (.A1(_01841_),
    .A2(\register_file[21][10] ),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14495_ (.A1(_02004_),
    .A2(_01840_),
    .A3(_02005_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14496_ (.A1(_01755_),
    .A2(\register_file[22][10] ),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14497_ (.A1(_01758_),
    .A2(\register_file[23][10] ),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14498_ (.A1(_02007_),
    .A2(_01757_),
    .A3(_02008_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14499_ (.A1(_02006_),
    .A2(_02009_),
    .A3(_01671_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14500_ (.A1(_02003_),
    .A2(_02010_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14501_ (.A1(_01993_),
    .A2(_02011_),
    .A3(_01930_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14502_ (.A1(_01932_),
    .A2(\register_file[8][10] ),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14503_ (.A1(_01676_),
    .A2(\register_file[9][10] ),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14504_ (.A1(_02013_),
    .A2(_02014_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14505_ (.A1(_02015_),
    .A2(_01853_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14506_ (.A1(_02016_),
    .A2(_01855_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14507_ (.A1(_01682_),
    .A2(\register_file[11][10] ),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14508_ (.A1(_01684_),
    .A2(\register_file[10][10] ),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14509_ (.A1(_02018_),
    .A2(_02019_),
    .B(_01859_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14510_ (.A1(_02017_),
    .A2(_02020_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14511_ (.A1(_01688_),
    .A2(\register_file[12][10] ),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14512_ (.A1(_01776_),
    .A2(\register_file[13][10] ),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14513_ (.A1(_02022_),
    .A2(_01775_),
    .A3(_02023_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14514_ (.I(_01161_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14515_ (.A1(_02025_),
    .A2(\register_file[14][10] ),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14516_ (.I(_01142_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14517_ (.A1(_02027_),
    .A2(\register_file[15][10] ),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14518_ (.A1(_02026_),
    .A2(_01694_),
    .A3(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14519_ (.I(_01147_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14520_ (.A1(_02024_),
    .A2(_02029_),
    .A3(_02030_),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14521_ (.A1(_02021_),
    .A2(_02031_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14522_ (.I(_01151_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14523_ (.A1(_02033_),
    .A2(\register_file[6][10] ),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14524_ (.I(\register_file[7][10] ),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14525_ (.A1(_02035_),
    .A2(_01786_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14526_ (.A1(_02034_),
    .A2(_02036_),
    .A3(_01702_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14527_ (.I(\register_file[4][10] ),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14528_ (.A1(_01954_),
    .A2(_02038_),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14529_ (.I(\register_file[5][10] ),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14530_ (.A1(_02040_),
    .A2(_01707_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14531_ (.A1(_02039_),
    .A2(_02041_),
    .A3(_01709_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14532_ (.A1(_02037_),
    .A2(_02042_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14533_ (.A1(_02043_),
    .A2(_01961_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14534_ (.I(_01176_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14535_ (.A1(_01713_),
    .A2(\register_file[2][10] ),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14536_ (.I(\register_file[3][10] ),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14537_ (.A1(_02047_),
    .A2(_01883_),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14538_ (.A1(_02045_),
    .A2(_02046_),
    .A3(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14539_ (.A1(_01800_),
    .A2(\register_file[1][10] ),
    .B(_01801_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14540_ (.A1(_02049_),
    .A2(_02050_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14541_ (.I(_02051_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14542_ (.A1(_02044_),
    .A2(_02052_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14543_ (.I(_01194_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14544_ (.A1(_02032_),
    .A2(_02053_),
    .A3(_02054_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14545_ (.I(_01200_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14546_ (.A1(_02012_),
    .A2(_02055_),
    .B(_02056_),
    .ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14547_ (.I(_00994_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14548_ (.A1(_02057_),
    .A2(\register_file[24][11] ),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14549_ (.A1(_01973_),
    .A2(\register_file[25][11] ),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14550_ (.A1(_02058_),
    .A2(_02059_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14551_ (.A1(_02060_),
    .A2(_01976_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14552_ (.A1(_02061_),
    .A2(_01811_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14553_ (.A1(_01813_),
    .A2(\register_file[27][11] ),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14554_ (.A1(_01980_),
    .A2(\register_file[26][11] ),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14555_ (.A1(_02063_),
    .A2(_02064_),
    .B(_01982_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14556_ (.A1(_02062_),
    .A2(_02065_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14557_ (.A1(_01818_),
    .A2(\register_file[28][11] ),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14558_ (.A1(_01986_),
    .A2(\register_file[29][11] ),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14559_ (.A1(_02067_),
    .A2(_01901_),
    .A3(_02068_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14560_ (.A1(_01904_),
    .A2(\register_file[30][11] ),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14561_ (.I(_01649_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14562_ (.A1(_02071_),
    .A2(\register_file[31][11] ),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14563_ (.A1(_02070_),
    .A2(_01906_),
    .A3(_02072_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14564_ (.A1(_02069_),
    .A2(_02073_),
    .A3(_01825_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14565_ (.A1(_02066_),
    .A2(_02074_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14566_ (.A1(_01994_),
    .A2(\register_file[16][11] ),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14567_ (.A1(_01741_),
    .A2(\register_file[17][11] ),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14568_ (.A1(_02076_),
    .A2(_02077_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14569_ (.A1(_02078_),
    .A2(_01914_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14570_ (.A1(_02079_),
    .A2(_01832_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14571_ (.A1(_01746_),
    .A2(\register_file[19][11] ),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14572_ (.A1(_01835_),
    .A2(\register_file[18][11] ),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14573_ (.A1(_02081_),
    .A2(_02082_),
    .B(_01919_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14574_ (.A1(_02080_),
    .A2(_02083_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14575_ (.A1(_01751_),
    .A2(\register_file[20][11] ),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14576_ (.A1(_01841_),
    .A2(\register_file[21][11] ),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14577_ (.A1(_02085_),
    .A2(_01840_),
    .A3(_02086_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14578_ (.A1(_01755_),
    .A2(\register_file[22][11] ),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14579_ (.A1(_01758_),
    .A2(\register_file[23][11] ),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14580_ (.A1(_02088_),
    .A2(_01757_),
    .A3(_02089_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14581_ (.I(_01670_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14582_ (.A1(_02087_),
    .A2(_02090_),
    .A3(_02091_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14583_ (.A1(_02084_),
    .A2(_02092_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14584_ (.A1(_02075_),
    .A2(_02093_),
    .A3(_01930_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14585_ (.A1(_01932_),
    .A2(\register_file[8][11] ),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14586_ (.I(_01110_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14587_ (.A1(_02096_),
    .A2(\register_file[9][11] ),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14588_ (.A1(_02095_),
    .A2(_02097_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14589_ (.A1(_02098_),
    .A2(_01853_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14590_ (.A1(_02099_),
    .A2(_01855_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14591_ (.I(_01681_),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14592_ (.A1(_02101_),
    .A2(\register_file[11][11] ),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14593_ (.I(_01122_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14594_ (.A1(_02103_),
    .A2(\register_file[10][11] ),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14595_ (.A1(_02102_),
    .A2(_02104_),
    .B(_01859_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14596_ (.A1(_02100_),
    .A2(_02105_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14597_ (.I(_01129_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14598_ (.A1(_02107_),
    .A2(\register_file[12][11] ),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14599_ (.A1(_01776_),
    .A2(\register_file[13][11] ),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14600_ (.A1(_02108_),
    .A2(_01775_),
    .A3(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14601_ (.A1(_02025_),
    .A2(\register_file[14][11] ),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14602_ (.I(_01693_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14603_ (.A1(_02027_),
    .A2(\register_file[15][11] ),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14604_ (.A1(_02111_),
    .A2(_02112_),
    .A3(_02113_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14605_ (.A1(_02110_),
    .A2(_02114_),
    .A3(_02030_),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14606_ (.A1(_02106_),
    .A2(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14607_ (.A1(_02033_),
    .A2(\register_file[6][11] ),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14608_ (.I(\register_file[7][11] ),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14609_ (.A1(_02118_),
    .A2(_01786_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14610_ (.I(_01158_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14611_ (.A1(_02117_),
    .A2(_02119_),
    .A3(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14612_ (.I(\register_file[4][11] ),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14613_ (.A1(_01954_),
    .A2(_02122_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14614_ (.I(\register_file[5][11] ),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14615_ (.I(_01166_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14616_ (.A1(_02124_),
    .A2(_02125_),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14617_ (.I(_01169_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14618_ (.A1(_02123_),
    .A2(_02126_),
    .A3(_02127_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14619_ (.A1(_02121_),
    .A2(_02128_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14620_ (.A1(_02129_),
    .A2(_01961_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14621_ (.I(_01277_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14622_ (.A1(_02131_),
    .A2(\register_file[2][11] ),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14623_ (.I(\register_file[3][11] ),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14624_ (.A1(_02133_),
    .A2(_01883_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14625_ (.A1(_02045_),
    .A2(_02132_),
    .A3(_02134_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14626_ (.A1(_01800_),
    .A2(\register_file[1][11] ),
    .B(_01801_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14627_ (.A1(_02135_),
    .A2(_02136_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14628_ (.I(_02137_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14629_ (.A1(_02130_),
    .A2(_02138_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14630_ (.A1(_02116_),
    .A2(_02139_),
    .A3(_02054_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14631_ (.A1(_02094_),
    .A2(_02140_),
    .B(_02056_),
    .ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14632_ (.A1(_02057_),
    .A2(\register_file[24][12] ),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14633_ (.A1(_01973_),
    .A2(\register_file[25][12] ),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14634_ (.A1(_02141_),
    .A2(_02142_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14635_ (.A1(_02143_),
    .A2(_01976_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14636_ (.A1(_02144_),
    .A2(_01811_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14637_ (.A1(_01813_),
    .A2(\register_file[27][12] ),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14638_ (.A1(_01980_),
    .A2(\register_file[26][12] ),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14639_ (.A1(_02146_),
    .A2(_02147_),
    .B(_01982_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14640_ (.A1(_02145_),
    .A2(_02148_),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14641_ (.A1(_01818_),
    .A2(\register_file[28][12] ),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14642_ (.A1(_01986_),
    .A2(\register_file[29][12] ),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14643_ (.A1(_02150_),
    .A2(_01901_),
    .A3(_02151_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14644_ (.A1(_01904_),
    .A2(\register_file[30][12] ),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14645_ (.A1(_02071_),
    .A2(\register_file[31][12] ),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14646_ (.A1(_02153_),
    .A2(_01906_),
    .A3(_02154_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14647_ (.A1(_02152_),
    .A2(_02155_),
    .A3(_01825_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14648_ (.A1(_02149_),
    .A2(_02156_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14649_ (.A1(_01994_),
    .A2(\register_file[16][12] ),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14650_ (.I(_01307_),
    .Z(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14651_ (.A1(_02159_),
    .A2(\register_file[17][12] ),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14652_ (.A1(_02158_),
    .A2(_02160_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14653_ (.A1(_02161_),
    .A2(_01914_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14654_ (.A1(_02162_),
    .A2(_01832_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14655_ (.I(_01119_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14656_ (.A1(_02164_),
    .A2(\register_file[19][12] ),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14657_ (.A1(_01835_),
    .A2(\register_file[18][12] ),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14658_ (.A1(_02165_),
    .A2(_02166_),
    .B(_01919_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14659_ (.A1(_02163_),
    .A2(_02167_),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14660_ (.I(_01318_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14661_ (.A1(_02169_),
    .A2(\register_file[20][12] ),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14662_ (.A1(_01841_),
    .A2(\register_file[21][12] ),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14663_ (.A1(_02170_),
    .A2(_01840_),
    .A3(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14664_ (.I(_01089_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14665_ (.A1(_02173_),
    .A2(\register_file[22][12] ),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14666_ (.I(_01325_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14667_ (.I(_01096_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14668_ (.A1(_02176_),
    .A2(\register_file[23][12] ),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14669_ (.A1(_02174_),
    .A2(_02175_),
    .A3(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14670_ (.A1(_02172_),
    .A2(_02178_),
    .A3(_02091_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14671_ (.A1(_02168_),
    .A2(_02179_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14672_ (.A1(_02157_),
    .A2(_02180_),
    .A3(_01930_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14673_ (.A1(_01932_),
    .A2(\register_file[8][12] ),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14674_ (.A1(_02096_),
    .A2(\register_file[9][12] ),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14675_ (.A1(_02182_),
    .A2(_02183_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14676_ (.A1(_02184_),
    .A2(_01853_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14677_ (.A1(_02185_),
    .A2(_01855_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14678_ (.A1(_02101_),
    .A2(\register_file[11][12] ),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14679_ (.A1(_02103_),
    .A2(\register_file[10][12] ),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14680_ (.A1(_02187_),
    .A2(_02188_),
    .B(_01859_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14681_ (.A1(_02186_),
    .A2(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14682_ (.A1(_02107_),
    .A2(\register_file[12][12] ),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14683_ (.I(_01774_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14684_ (.I(_01047_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14685_ (.A1(_02193_),
    .A2(\register_file[13][12] ),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14686_ (.A1(_02191_),
    .A2(_02192_),
    .A3(_02194_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14687_ (.A1(_02025_),
    .A2(\register_file[14][12] ),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14688_ (.A1(_02027_),
    .A2(\register_file[15][12] ),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14689_ (.A1(_02196_),
    .A2(_02112_),
    .A3(_02197_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14690_ (.A1(_02195_),
    .A2(_02198_),
    .A3(_02030_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14691_ (.A1(_02190_),
    .A2(_02199_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14692_ (.A1(_02033_),
    .A2(\register_file[6][12] ),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14693_ (.I(\register_file[7][12] ),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14694_ (.I(_01354_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14695_ (.A1(_02202_),
    .A2(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14696_ (.A1(_02201_),
    .A2(_02204_),
    .A3(_02120_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14697_ (.I(\register_file[4][12] ),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14698_ (.A1(_01954_),
    .A2(_02206_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14699_ (.I(\register_file[5][12] ),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14700_ (.A1(_02208_),
    .A2(_02125_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14701_ (.A1(_02207_),
    .A2(_02209_),
    .A3(_02127_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14702_ (.A1(_02205_),
    .A2(_02210_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14703_ (.A1(_02211_),
    .A2(_01961_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14704_ (.A1(_02131_),
    .A2(\register_file[2][12] ),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14705_ (.I(\register_file[3][12] ),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14706_ (.A1(_02214_),
    .A2(_01883_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14707_ (.A1(_02045_),
    .A2(_02213_),
    .A3(_02215_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14708_ (.I(_01185_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14709_ (.I(_01370_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14710_ (.A1(_02217_),
    .A2(\register_file[1][12] ),
    .B(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14711_ (.A1(_02216_),
    .A2(_02219_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14712_ (.I(_02220_),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14713_ (.A1(_02212_),
    .A2(_02221_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14714_ (.A1(_02200_),
    .A2(_02222_),
    .A3(_02054_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14715_ (.A1(_02181_),
    .A2(_02223_),
    .B(_02056_),
    .ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14716_ (.A1(_02057_),
    .A2(\register_file[24][13] ),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14717_ (.A1(_01973_),
    .A2(\register_file[25][13] ),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14718_ (.A1(_02224_),
    .A2(_02225_),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14719_ (.A1(_02226_),
    .A2(_01976_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14720_ (.I(_01065_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14721_ (.A1(_02227_),
    .A2(_02228_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14722_ (.I(_01014_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14723_ (.A1(_02230_),
    .A2(\register_file[27][13] ),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14724_ (.A1(_01980_),
    .A2(\register_file[26][13] ),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14725_ (.A1(_02231_),
    .A2(_02232_),
    .B(_01982_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14726_ (.A1(_02229_),
    .A2(_02233_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14727_ (.I(_01080_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14728_ (.A1(_02235_),
    .A2(\register_file[28][13] ),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14729_ (.A1(_01986_),
    .A2(\register_file[29][13] ),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14730_ (.A1(_02236_),
    .A2(_01901_),
    .A3(_02237_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14731_ (.A1(_01904_),
    .A2(\register_file[30][13] ),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14732_ (.A1(_02071_),
    .A2(\register_file[31][13] ),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14733_ (.A1(_02239_),
    .A2(_01906_),
    .A3(_02240_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14734_ (.I(_01100_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14735_ (.A1(_02238_),
    .A2(_02241_),
    .A3(_02242_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14736_ (.A1(_02234_),
    .A2(_02243_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14737_ (.A1(_01994_),
    .A2(\register_file[16][13] ),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14738_ (.A1(_02159_),
    .A2(\register_file[17][13] ),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14739_ (.A1(_02245_),
    .A2(_02246_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14740_ (.A1(_02247_),
    .A2(_01914_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14741_ (.I(_01008_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14742_ (.A1(_02248_),
    .A2(_02249_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14743_ (.A1(_02164_),
    .A2(\register_file[19][13] ),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14744_ (.I(_01404_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14745_ (.A1(_02252_),
    .A2(\register_file[18][13] ),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14746_ (.A1(_02251_),
    .A2(_02253_),
    .B(_01919_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14747_ (.A1(_02250_),
    .A2(_02254_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14748_ (.A1(_02169_),
    .A2(\register_file[20][13] ),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14749_ (.I(_01132_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14750_ (.I(_01085_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14751_ (.A1(_02258_),
    .A2(\register_file[21][13] ),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14752_ (.A1(_02256_),
    .A2(_02257_),
    .A3(_02259_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14753_ (.A1(_02173_),
    .A2(\register_file[22][13] ),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14754_ (.A1(_02176_),
    .A2(\register_file[23][13] ),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14755_ (.A1(_02261_),
    .A2(_02175_),
    .A3(_02262_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14756_ (.A1(_02260_),
    .A2(_02263_),
    .A3(_02091_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14757_ (.A1(_02255_),
    .A2(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14758_ (.A1(_02244_),
    .A2(_02265_),
    .A3(_01930_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14759_ (.A1(_01932_),
    .A2(\register_file[8][13] ),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14760_ (.A1(_02096_),
    .A2(\register_file[9][13] ),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14761_ (.A1(_02267_),
    .A2(_02268_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14762_ (.I(_01423_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14763_ (.A1(_02269_),
    .A2(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14764_ (.I(_01426_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14765_ (.A1(_02271_),
    .A2(_02272_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14766_ (.A1(_02101_),
    .A2(\register_file[11][13] ),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14767_ (.A1(_02103_),
    .A2(\register_file[10][13] ),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14768_ (.I(_01125_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14769_ (.A1(_02274_),
    .A2(_02275_),
    .B(_02276_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14770_ (.A1(_02273_),
    .A2(_02277_),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14771_ (.A1(_02107_),
    .A2(\register_file[12][13] ),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14772_ (.A1(_02193_),
    .A2(\register_file[13][13] ),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14773_ (.A1(_02279_),
    .A2(_02192_),
    .A3(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14774_ (.A1(_02025_),
    .A2(\register_file[14][13] ),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14775_ (.A1(_02027_),
    .A2(\register_file[15][13] ),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14776_ (.A1(_02282_),
    .A2(_02112_),
    .A3(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14777_ (.A1(_02281_),
    .A2(_02284_),
    .A3(_02030_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14778_ (.A1(_02278_),
    .A2(_02285_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14779_ (.A1(_02033_),
    .A2(\register_file[6][13] ),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14780_ (.I(\register_file[7][13] ),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14781_ (.A1(_02288_),
    .A2(_02203_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14782_ (.A1(_02287_),
    .A2(_02289_),
    .A3(_02120_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14783_ (.I(\register_file[4][13] ),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14784_ (.A1(_01954_),
    .A2(_02291_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14785_ (.I(\register_file[5][13] ),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14786_ (.A1(_02293_),
    .A2(_02125_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14787_ (.A1(_02292_),
    .A2(_02294_),
    .A3(_02127_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14788_ (.A1(_02290_),
    .A2(_02295_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14789_ (.A1(_02296_),
    .A2(_01961_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14790_ (.A1(_02131_),
    .A2(\register_file[2][13] ),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14791_ (.I(\register_file[3][13] ),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14792_ (.I(_01155_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14793_ (.A1(_02299_),
    .A2(_02300_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14794_ (.A1(_02045_),
    .A2(_02298_),
    .A3(_02301_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14795_ (.A1(_02217_),
    .A2(\register_file[1][13] ),
    .B(_02218_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14796_ (.A1(_02302_),
    .A2(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14797_ (.I(_02304_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14798_ (.A1(_02297_),
    .A2(_02305_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14799_ (.A1(_02286_),
    .A2(_02306_),
    .A3(_02054_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14800_ (.A1(_02266_),
    .A2(_02307_),
    .B(_02056_),
    .ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14801_ (.A1(_02057_),
    .A2(\register_file[24][14] ),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14802_ (.A1(_01973_),
    .A2(\register_file[25][14] ),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14803_ (.A1(_02308_),
    .A2(_02309_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14804_ (.A1(_02310_),
    .A2(_01976_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14805_ (.A1(_02311_),
    .A2(_02228_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14806_ (.A1(_02230_),
    .A2(\register_file[27][14] ),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14807_ (.A1(_01980_),
    .A2(\register_file[26][14] ),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14808_ (.A1(_02313_),
    .A2(_02314_),
    .B(_01982_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14809_ (.A1(_02312_),
    .A2(_02315_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14810_ (.A1(_02235_),
    .A2(\register_file[28][14] ),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14811_ (.I(_01035_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14812_ (.A1(_01986_),
    .A2(\register_file[29][14] ),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14813_ (.A1(_02317_),
    .A2(_02318_),
    .A3(_02319_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14814_ (.I(_01071_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14815_ (.A1(_02321_),
    .A2(\register_file[30][14] ),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14816_ (.I(_01045_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14817_ (.A1(_02071_),
    .A2(\register_file[31][14] ),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14818_ (.A1(_02322_),
    .A2(_02323_),
    .A3(_02324_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14819_ (.A1(_02320_),
    .A2(_02325_),
    .A3(_02242_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14820_ (.A1(_02316_),
    .A2(_02326_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14821_ (.A1(_01994_),
    .A2(\register_file[16][14] ),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14822_ (.A1(_02159_),
    .A2(\register_file[17][14] ),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14823_ (.A1(_02328_),
    .A2(_02329_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14824_ (.I(_01114_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14825_ (.A1(_02330_),
    .A2(_02331_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14826_ (.A1(_02332_),
    .A2(_02249_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14827_ (.A1(_02164_),
    .A2(\register_file[19][14] ),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14828_ (.A1(_02252_),
    .A2(\register_file[18][14] ),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14829_ (.I(_01075_),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14830_ (.A1(_02334_),
    .A2(_02335_),
    .B(_02336_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14831_ (.A1(_02333_),
    .A2(_02337_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14832_ (.A1(_02169_),
    .A2(\register_file[20][14] ),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14833_ (.A1(_02258_),
    .A2(\register_file[21][14] ),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14834_ (.A1(_02339_),
    .A2(_02257_),
    .A3(_02340_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14835_ (.A1(_02173_),
    .A2(\register_file[22][14] ),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14836_ (.A1(_02176_),
    .A2(\register_file[23][14] ),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14837_ (.A1(_02342_),
    .A2(_02175_),
    .A3(_02343_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14838_ (.A1(_02341_),
    .A2(_02344_),
    .A3(_02091_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14839_ (.A1(_02338_),
    .A2(_02345_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14840_ (.I(_01104_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14841_ (.A1(_02327_),
    .A2(_02346_),
    .A3(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14842_ (.I(_01079_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14843_ (.A1(_02349_),
    .A2(\register_file[8][14] ),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14844_ (.A1(_02096_),
    .A2(\register_file[9][14] ),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14845_ (.A1(_02350_),
    .A2(_02351_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14846_ (.A1(_02352_),
    .A2(_02270_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14847_ (.A1(_02353_),
    .A2(_02272_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14848_ (.A1(_02101_),
    .A2(\register_file[11][14] ),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14849_ (.A1(_02103_),
    .A2(\register_file[10][14] ),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14850_ (.A1(_02355_),
    .A2(_02356_),
    .B(_02276_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14851_ (.A1(_02354_),
    .A2(_02357_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14852_ (.A1(_02107_),
    .A2(\register_file[12][14] ),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14853_ (.A1(_02193_),
    .A2(\register_file[13][14] ),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14854_ (.A1(_02359_),
    .A2(_02192_),
    .A3(_02360_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14855_ (.A1(_02025_),
    .A2(\register_file[14][14] ),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14856_ (.A1(_02027_),
    .A2(\register_file[15][14] ),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14857_ (.A1(_02362_),
    .A2(_02112_),
    .A3(_02363_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14858_ (.A1(_02361_),
    .A2(_02364_),
    .A3(_02030_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14859_ (.A1(_02358_),
    .A2(_02365_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14860_ (.A1(_02033_),
    .A2(\register_file[6][14] ),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14861_ (.I(\register_file[7][14] ),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14862_ (.A1(_02368_),
    .A2(_02203_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14863_ (.A1(_02367_),
    .A2(_02369_),
    .A3(_02120_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14864_ (.I(_01530_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14865_ (.I(\register_file[4][14] ),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14866_ (.A1(_02371_),
    .A2(_02372_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14867_ (.I(\register_file[5][14] ),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14868_ (.A1(_02374_),
    .A2(_02125_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14869_ (.A1(_02373_),
    .A2(_02375_),
    .A3(_02127_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14870_ (.A1(_02370_),
    .A2(_02376_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14871_ (.I(_01146_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14872_ (.A1(_02377_),
    .A2(_02378_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14873_ (.A1(_02131_),
    .A2(\register_file[2][14] ),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14874_ (.I(\register_file[3][14] ),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14875_ (.A1(_02381_),
    .A2(_02300_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14876_ (.A1(_02045_),
    .A2(_02380_),
    .A3(_02382_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14877_ (.A1(_02217_),
    .A2(\register_file[1][14] ),
    .B(_02218_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14878_ (.A1(_02383_),
    .A2(_02384_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14879_ (.I(_02385_),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14880_ (.A1(_02379_),
    .A2(_02386_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14881_ (.A1(_02366_),
    .A2(_02387_),
    .A3(_02054_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14882_ (.A1(_02348_),
    .A2(_02388_),
    .B(_02056_),
    .ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14883_ (.A1(_02057_),
    .A2(\register_file[24][15] ),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14884_ (.I(_01058_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14885_ (.A1(_02390_),
    .A2(\register_file[25][15] ),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14886_ (.A1(_02389_),
    .A2(_02391_),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14887_ (.I(_01062_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14888_ (.A1(_02392_),
    .A2(_02393_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14889_ (.A1(_02394_),
    .A2(_02228_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14890_ (.A1(_02230_),
    .A2(\register_file[27][15] ),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14891_ (.I(_01042_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14892_ (.A1(_02397_),
    .A2(\register_file[26][15] ),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14893_ (.I(_01559_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14894_ (.A1(_02396_),
    .A2(_02398_),
    .B(_02399_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14895_ (.A1(_02395_),
    .A2(_02400_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14896_ (.A1(_02235_),
    .A2(\register_file[28][15] ),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14897_ (.I(_01038_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14898_ (.A1(_02403_),
    .A2(\register_file[29][15] ),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14899_ (.A1(_02402_),
    .A2(_02318_),
    .A3(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14900_ (.A1(_02321_),
    .A2(\register_file[30][15] ),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14901_ (.A1(_02071_),
    .A2(\register_file[31][15] ),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14902_ (.A1(_02406_),
    .A2(_02323_),
    .A3(_02407_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14903_ (.A1(_02405_),
    .A2(_02408_),
    .A3(_02242_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14904_ (.A1(_02401_),
    .A2(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14905_ (.I(_01107_),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14906_ (.A1(_02411_),
    .A2(\register_file[16][15] ),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14907_ (.A1(_02159_),
    .A2(\register_file[17][15] ),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14908_ (.A1(_02412_),
    .A2(_02413_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14909_ (.A1(_02414_),
    .A2(_02331_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14910_ (.A1(_02415_),
    .A2(_02249_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14911_ (.A1(_02164_),
    .A2(\register_file[19][15] ),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14912_ (.A1(_02252_),
    .A2(\register_file[18][15] ),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14913_ (.A1(_02417_),
    .A2(_02418_),
    .B(_02336_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14914_ (.A1(_02416_),
    .A2(_02419_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14915_ (.A1(_02169_),
    .A2(\register_file[20][15] ),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14916_ (.A1(_02258_),
    .A2(\register_file[21][15] ),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14917_ (.A1(_02421_),
    .A2(_02257_),
    .A3(_02422_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14918_ (.A1(_02173_),
    .A2(\register_file[22][15] ),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14919_ (.A1(_02176_),
    .A2(\register_file[23][15] ),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14920_ (.A1(_02424_),
    .A2(_02175_),
    .A3(_02425_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14921_ (.A1(_02423_),
    .A2(_02426_),
    .A3(_02091_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14922_ (.A1(_02420_),
    .A2(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14923_ (.A1(_02410_),
    .A2(_02428_),
    .A3(_02347_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14924_ (.A1(_02349_),
    .A2(\register_file[8][15] ),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14925_ (.A1(_02096_),
    .A2(\register_file[9][15] ),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14926_ (.A1(_02430_),
    .A2(_02431_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14927_ (.A1(_02432_),
    .A2(_02270_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14928_ (.A1(_02433_),
    .A2(_02272_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14929_ (.A1(_02101_),
    .A2(\register_file[11][15] ),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14930_ (.A1(_02103_),
    .A2(\register_file[10][15] ),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14931_ (.A1(_02435_),
    .A2(_02436_),
    .B(_02276_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14932_ (.A1(_02434_),
    .A2(_02437_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14933_ (.A1(_02107_),
    .A2(\register_file[12][15] ),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14934_ (.A1(_02193_),
    .A2(\register_file[13][15] ),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14935_ (.A1(_02439_),
    .A2(_02192_),
    .A3(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14936_ (.I(_01161_),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14937_ (.A1(_02442_),
    .A2(\register_file[14][15] ),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14938_ (.I(_01455_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14939_ (.A1(_02444_),
    .A2(\register_file[15][15] ),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14940_ (.A1(_02443_),
    .A2(_02112_),
    .A3(_02445_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14941_ (.I(_01147_),
    .Z(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14942_ (.A1(_02441_),
    .A2(_02446_),
    .A3(_02447_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14943_ (.A1(_02438_),
    .A2(_02448_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14944_ (.I(_01178_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14945_ (.A1(_02450_),
    .A2(\register_file[6][15] ),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14946_ (.I(\register_file[7][15] ),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14947_ (.A1(_02452_),
    .A2(_02203_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14948_ (.A1(_02451_),
    .A2(_02453_),
    .A3(_02120_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14949_ (.I(\register_file[4][15] ),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14950_ (.A1(_02371_),
    .A2(_02455_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14951_ (.I(\register_file[5][15] ),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14952_ (.A1(_02457_),
    .A2(_02125_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14953_ (.A1(_02456_),
    .A2(_02458_),
    .A3(_02127_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14954_ (.A1(_02454_),
    .A2(_02459_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14955_ (.A1(_02460_),
    .A2(_02378_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14956_ (.I(_01176_),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14957_ (.A1(_02131_),
    .A2(\register_file[2][15] ),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14958_ (.I(\register_file[3][15] ),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14959_ (.A1(_02464_),
    .A2(_02300_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14960_ (.A1(_02462_),
    .A2(_02463_),
    .A3(_02465_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14961_ (.A1(_02217_),
    .A2(\register_file[1][15] ),
    .B(_02218_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14962_ (.A1(_02466_),
    .A2(_02467_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14963_ (.I(_02468_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14964_ (.A1(_02461_),
    .A2(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14965_ (.I(_01194_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14966_ (.A1(_02449_),
    .A2(_02470_),
    .A3(_02471_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14967_ (.I(_01200_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14968_ (.A1(_02429_),
    .A2(_02472_),
    .B(_02473_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14969_ (.I(_00994_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14970_ (.A1(_02474_),
    .A2(\register_file[24][16] ),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14971_ (.A1(_02390_),
    .A2(\register_file[25][16] ),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14972_ (.A1(_02475_),
    .A2(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14973_ (.A1(_02477_),
    .A2(_02393_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14974_ (.A1(_02478_),
    .A2(_02228_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14975_ (.A1(_02230_),
    .A2(\register_file[27][16] ),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14976_ (.A1(_02397_),
    .A2(\register_file[26][16] ),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14977_ (.A1(_02480_),
    .A2(_02481_),
    .B(_02399_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14978_ (.A1(_02479_),
    .A2(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14979_ (.A1(_02235_),
    .A2(\register_file[28][16] ),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14980_ (.A1(_02403_),
    .A2(\register_file[29][16] ),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14981_ (.A1(_02484_),
    .A2(_02318_),
    .A3(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14982_ (.A1(_02321_),
    .A2(\register_file[30][16] ),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14983_ (.I(_01649_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14984_ (.A1(_02488_),
    .A2(\register_file[31][16] ),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14985_ (.A1(_02487_),
    .A2(_02323_),
    .A3(_02489_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14986_ (.A1(_02486_),
    .A2(_02490_),
    .A3(_02242_),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14987_ (.A1(_02483_),
    .A2(_02491_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14988_ (.A1(_02411_),
    .A2(\register_file[16][16] ),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14989_ (.A1(_02159_),
    .A2(\register_file[17][16] ),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14990_ (.A1(_02493_),
    .A2(_02494_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14991_ (.A1(_02495_),
    .A2(_02331_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14992_ (.A1(_02496_),
    .A2(_02249_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14993_ (.A1(_02164_),
    .A2(\register_file[19][16] ),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14994_ (.A1(_02252_),
    .A2(\register_file[18][16] ),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14995_ (.A1(_02498_),
    .A2(_02499_),
    .B(_02336_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14996_ (.A1(_02497_),
    .A2(_02500_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14997_ (.A1(_02169_),
    .A2(\register_file[20][16] ),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14998_ (.A1(_02258_),
    .A2(\register_file[21][16] ),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14999_ (.A1(_02502_),
    .A2(_02257_),
    .A3(_02503_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15000_ (.A1(_02173_),
    .A2(\register_file[22][16] ),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15001_ (.A1(_02176_),
    .A2(\register_file[23][16] ),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15002_ (.A1(_02505_),
    .A2(_02175_),
    .A3(_02506_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15003_ (.I(_01670_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15004_ (.A1(_02504_),
    .A2(_02507_),
    .A3(_02508_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15005_ (.A1(_02501_),
    .A2(_02509_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15006_ (.A1(_02492_),
    .A2(_02510_),
    .A3(_02347_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15007_ (.A1(_02349_),
    .A2(\register_file[8][16] ),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15008_ (.I(_01110_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15009_ (.A1(_02513_),
    .A2(\register_file[9][16] ),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15010_ (.A1(_02512_),
    .A2(_02514_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15011_ (.A1(_02515_),
    .A2(_02270_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15012_ (.A1(_02516_),
    .A2(_02272_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15013_ (.I(_01681_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15014_ (.A1(_02518_),
    .A2(\register_file[11][16] ),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15015_ (.I(_01138_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15016_ (.A1(_02520_),
    .A2(\register_file[10][16] ),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15017_ (.A1(_02519_),
    .A2(_02521_),
    .B(_02276_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15018_ (.A1(_02517_),
    .A2(_02522_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15019_ (.I(_01129_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15020_ (.A1(_02524_),
    .A2(\register_file[12][16] ),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15021_ (.A1(_02193_),
    .A2(\register_file[13][16] ),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15022_ (.A1(_02525_),
    .A2(_02192_),
    .A3(_02526_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15023_ (.A1(_02442_),
    .A2(\register_file[14][16] ),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15024_ (.I(_01693_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15025_ (.A1(_02444_),
    .A2(\register_file[15][16] ),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15026_ (.A1(_02528_),
    .A2(_02529_),
    .A3(_02530_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15027_ (.A1(_02527_),
    .A2(_02531_),
    .A3(_02447_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15028_ (.A1(_02523_),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15029_ (.A1(_02450_),
    .A2(\register_file[6][16] ),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15030_ (.I(\register_file[7][16] ),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15031_ (.A1(_02535_),
    .A2(_02203_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15032_ (.I(_01158_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15033_ (.A1(_02534_),
    .A2(_02536_),
    .A3(_02537_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15034_ (.I(\register_file[4][16] ),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15035_ (.A1(_02371_),
    .A2(_02539_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15036_ (.I(\register_file[5][16] ),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15037_ (.I(_01166_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15038_ (.A1(_02541_),
    .A2(_02542_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15039_ (.I(_01169_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15040_ (.A1(_02540_),
    .A2(_02543_),
    .A3(_02544_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15041_ (.A1(_02538_),
    .A2(_02545_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15042_ (.A1(_02546_),
    .A2(_02378_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15043_ (.I(_01277_),
    .Z(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15044_ (.A1(_02548_),
    .A2(\register_file[2][16] ),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15045_ (.I(\register_file[3][16] ),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15046_ (.A1(_02550_),
    .A2(_02300_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15047_ (.A1(_02462_),
    .A2(_02549_),
    .A3(_02551_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15048_ (.A1(_02217_),
    .A2(\register_file[1][16] ),
    .B(_02218_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15049_ (.A1(_02552_),
    .A2(_02553_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15050_ (.I(_02554_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15051_ (.A1(_02547_),
    .A2(_02555_),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15052_ (.A1(_02533_),
    .A2(_02556_),
    .A3(_02471_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15053_ (.A1(_02511_),
    .A2(_02557_),
    .B(_02473_),
    .ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15054_ (.A1(_02474_),
    .A2(\register_file[24][17] ),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15055_ (.A1(_02390_),
    .A2(\register_file[25][17] ),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15056_ (.A1(_02558_),
    .A2(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15057_ (.A1(_02560_),
    .A2(_02393_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15058_ (.A1(_02561_),
    .A2(_02228_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15059_ (.A1(_02230_),
    .A2(\register_file[27][17] ),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15060_ (.A1(_02397_),
    .A2(\register_file[26][17] ),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15061_ (.A1(_02563_),
    .A2(_02564_),
    .B(_02399_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15062_ (.A1(_02562_),
    .A2(_02565_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15063_ (.A1(_02235_),
    .A2(\register_file[28][17] ),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15064_ (.A1(_02403_),
    .A2(\register_file[29][17] ),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15065_ (.A1(_02567_),
    .A2(_02318_),
    .A3(_02568_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15066_ (.A1(_02321_),
    .A2(\register_file[30][17] ),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15067_ (.A1(_02488_),
    .A2(\register_file[31][17] ),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15068_ (.A1(_02570_),
    .A2(_02323_),
    .A3(_02571_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15069_ (.A1(_02569_),
    .A2(_02572_),
    .A3(_02242_),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15070_ (.A1(_02566_),
    .A2(_02573_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15071_ (.A1(_02411_),
    .A2(\register_file[16][17] ),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15072_ (.I(_01307_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15073_ (.A1(_02576_),
    .A2(\register_file[17][17] ),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15074_ (.A1(_02575_),
    .A2(_02577_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15075_ (.A1(_02578_),
    .A2(_02331_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15076_ (.A1(_02579_),
    .A2(_02249_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15077_ (.I(_01119_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15078_ (.A1(_02581_),
    .A2(\register_file[19][17] ),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15079_ (.A1(_02252_),
    .A2(\register_file[18][17] ),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15080_ (.A1(_02582_),
    .A2(_02583_),
    .B(_02336_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15081_ (.A1(_02580_),
    .A2(_02584_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15082_ (.I(_01318_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15083_ (.A1(_02586_),
    .A2(\register_file[20][17] ),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15084_ (.A1(_02258_),
    .A2(\register_file[21][17] ),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15085_ (.A1(_02587_),
    .A2(_02257_),
    .A3(_02588_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15086_ (.I(_01089_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15087_ (.A1(_02590_),
    .A2(\register_file[22][17] ),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15088_ (.I(_01093_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15089_ (.I(_01142_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15090_ (.A1(_02593_),
    .A2(\register_file[23][17] ),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15091_ (.A1(_02591_),
    .A2(_02592_),
    .A3(_02594_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15092_ (.A1(_02589_),
    .A2(_02595_),
    .A3(_02508_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15093_ (.A1(_02585_),
    .A2(_02596_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15094_ (.A1(_02574_),
    .A2(_02597_),
    .A3(_02347_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15095_ (.A1(_02349_),
    .A2(\register_file[8][17] ),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15096_ (.A1(_02513_),
    .A2(\register_file[9][17] ),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15097_ (.A1(_02599_),
    .A2(_02600_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15098_ (.A1(_02601_),
    .A2(_02270_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15099_ (.A1(_02602_),
    .A2(_02272_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15100_ (.A1(_02518_),
    .A2(\register_file[11][17] ),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15101_ (.A1(_02520_),
    .A2(\register_file[10][17] ),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15102_ (.A1(_02604_),
    .A2(_02605_),
    .B(_02276_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15103_ (.A1(_02603_),
    .A2(_02606_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15104_ (.A1(_02524_),
    .A2(\register_file[12][17] ),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15105_ (.I(_01774_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15106_ (.I(_01047_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15107_ (.A1(_02610_),
    .A2(\register_file[13][17] ),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15108_ (.A1(_02608_),
    .A2(_02609_),
    .A3(_02611_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15109_ (.A1(_02442_),
    .A2(\register_file[14][17] ),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15110_ (.A1(_02444_),
    .A2(\register_file[15][17] ),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15111_ (.A1(_02613_),
    .A2(_02529_),
    .A3(_02614_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15112_ (.A1(_02612_),
    .A2(_02615_),
    .A3(_02447_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15113_ (.A1(_02607_),
    .A2(_02616_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15114_ (.A1(_02450_),
    .A2(\register_file[6][17] ),
    .Z(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15115_ (.I(\register_file[7][17] ),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15116_ (.I(_01354_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15117_ (.A1(_02619_),
    .A2(_02620_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15118_ (.A1(_02618_),
    .A2(_02621_),
    .A3(_02537_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15119_ (.I(\register_file[4][17] ),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15120_ (.A1(_02371_),
    .A2(_02623_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15121_ (.I(\register_file[5][17] ),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15122_ (.A1(_02625_),
    .A2(_02542_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15123_ (.A1(_02624_),
    .A2(_02626_),
    .A3(_02544_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15124_ (.A1(_02622_),
    .A2(_02627_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15125_ (.A1(_02628_),
    .A2(_02378_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15126_ (.A1(_02548_),
    .A2(\register_file[2][17] ),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15127_ (.I(\register_file[3][17] ),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15128_ (.A1(_02631_),
    .A2(_02300_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15129_ (.A1(_02462_),
    .A2(_02630_),
    .A3(_02632_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15130_ (.I(_01185_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15131_ (.I(_01370_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15132_ (.A1(_02634_),
    .A2(\register_file[1][17] ),
    .B(_02635_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15133_ (.A1(_02633_),
    .A2(_02636_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15134_ (.I(_02637_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15135_ (.A1(_02629_),
    .A2(_02638_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15136_ (.A1(_02617_),
    .A2(_02639_),
    .A3(_02471_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15137_ (.A1(_02598_),
    .A2(_02640_),
    .B(_02473_),
    .ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15138_ (.A1(_02474_),
    .A2(\register_file[16][18] ),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15139_ (.A1(_02390_),
    .A2(\register_file[17][18] ),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15140_ (.A1(_02641_),
    .A2(_02642_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15141_ (.A1(_02643_),
    .A2(_02393_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15142_ (.A1(_02644_),
    .A2(_01292_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15143_ (.I(_01068_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15144_ (.A1(_02646_),
    .A2(\register_file[19][18] ),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15145_ (.A1(_02397_),
    .A2(\register_file[18][18] ),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15146_ (.A1(_02647_),
    .A2(_02648_),
    .B(_02399_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15147_ (.A1(_02645_),
    .A2(_02649_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15148_ (.I(_01080_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15149_ (.A1(_02651_),
    .A2(\register_file[20][18] ),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15150_ (.A1(_02403_),
    .A2(\register_file[21][18] ),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15151_ (.A1(_02652_),
    .A2(_02318_),
    .A3(_02653_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15152_ (.A1(_02321_),
    .A2(\register_file[22][18] ),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15153_ (.A1(_02488_),
    .A2(\register_file[23][18] ),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15154_ (.A1(_02655_),
    .A2(_02323_),
    .A3(_02656_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15155_ (.I(_01100_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15156_ (.A1(_02654_),
    .A2(_02657_),
    .A3(_02658_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15157_ (.A1(_02650_),
    .A2(_02659_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15158_ (.A1(_02411_),
    .A2(\register_file[24][18] ),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15159_ (.A1(_02576_),
    .A2(\register_file[25][18] ),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15160_ (.A1(_02661_),
    .A2(_02662_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15161_ (.A1(_02663_),
    .A2(_02331_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15162_ (.A1(_02664_),
    .A2(_01225_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15163_ (.A1(_02581_),
    .A2(\register_file[27][18] ),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15164_ (.I(_01404_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15165_ (.A1(_02667_),
    .A2(\register_file[26][18] ),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15166_ (.A1(_02666_),
    .A2(_02668_),
    .B(_02336_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15167_ (.A1(_02665_),
    .A2(_02669_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15168_ (.A1(_02586_),
    .A2(\register_file[28][18] ),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15169_ (.I(_01132_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15170_ (.I(_01134_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15171_ (.A1(_02673_),
    .A2(\register_file[29][18] ),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15172_ (.A1(_02671_),
    .A2(_02672_),
    .A3(_02674_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15173_ (.A1(_02590_),
    .A2(\register_file[30][18] ),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15174_ (.A1(_02593_),
    .A2(\register_file[31][18] ),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15175_ (.A1(_02676_),
    .A2(_02592_),
    .A3(_02677_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15176_ (.A1(_02675_),
    .A2(_02678_),
    .A3(_02508_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15177_ (.A1(_02670_),
    .A2(_02679_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15178_ (.A1(_02660_),
    .A2(_02680_),
    .A3(_02347_),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15179_ (.A1(_02349_),
    .A2(\register_file[8][18] ),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15180_ (.A1(_02513_),
    .A2(\register_file[9][18] ),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15181_ (.A1(_02682_),
    .A2(_02683_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15182_ (.I(_01423_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15183_ (.A1(_02684_),
    .A2(_02685_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15184_ (.I(_01426_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15185_ (.A1(_02686_),
    .A2(_02687_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15186_ (.A1(_02518_),
    .A2(\register_file[11][18] ),
    .ZN(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15187_ (.A1(_02520_),
    .A2(\register_file[10][18] ),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15188_ (.I(_01074_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15189_ (.A1(_02689_),
    .A2(_02690_),
    .B(_02691_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15190_ (.A1(_02688_),
    .A2(_02692_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15191_ (.A1(_02524_),
    .A2(\register_file[12][18] ),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15192_ (.A1(_02610_),
    .A2(\register_file[13][18] ),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15193_ (.A1(_02694_),
    .A2(_02609_),
    .A3(_02695_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15194_ (.A1(_02442_),
    .A2(\register_file[14][18] ),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15195_ (.A1(_02444_),
    .A2(\register_file[15][18] ),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15196_ (.A1(_02697_),
    .A2(_02529_),
    .A3(_02698_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15197_ (.A1(_02696_),
    .A2(_02699_),
    .A3(_02447_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15198_ (.A1(_02693_),
    .A2(_02700_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15199_ (.A1(_02450_),
    .A2(\register_file[6][18] ),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15200_ (.I(\register_file[7][18] ),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15201_ (.A1(_02703_),
    .A2(_02620_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15202_ (.A1(_02702_),
    .A2(_02704_),
    .A3(_02537_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15203_ (.I(\register_file[4][18] ),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15204_ (.A1(_02371_),
    .A2(_02706_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15205_ (.I(\register_file[5][18] ),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15206_ (.A1(_02708_),
    .A2(_02542_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15207_ (.A1(_02707_),
    .A2(_02709_),
    .A3(_02544_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15208_ (.A1(_02705_),
    .A2(_02710_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15209_ (.A1(_02711_),
    .A2(_02378_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15210_ (.A1(_02548_),
    .A2(\register_file[2][18] ),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15211_ (.I(\register_file[3][18] ),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15212_ (.I(_01155_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15213_ (.A1(_02714_),
    .A2(_02715_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15214_ (.A1(_02462_),
    .A2(_02713_),
    .A3(_02716_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15215_ (.A1(_02634_),
    .A2(\register_file[1][18] ),
    .B(_02635_),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15216_ (.A1(_02717_),
    .A2(_02718_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15217_ (.I(_02719_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15218_ (.A1(_02712_),
    .A2(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15219_ (.A1(_02701_),
    .A2(_02721_),
    .A3(_02471_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15220_ (.A1(_02681_),
    .A2(_02722_),
    .B(_02473_),
    .ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15221_ (.A1(_02474_),
    .A2(\register_file[16][19] ),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15222_ (.A1(_02390_),
    .A2(\register_file[17][19] ),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15223_ (.A1(_02723_),
    .A2(_02724_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15224_ (.A1(_02725_),
    .A2(_02393_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15225_ (.A1(_02726_),
    .A2(_01292_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15226_ (.A1(_02646_),
    .A2(\register_file[19][19] ),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15227_ (.A1(_02397_),
    .A2(\register_file[18][19] ),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15228_ (.A1(_02728_),
    .A2(_02729_),
    .B(_02399_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15229_ (.A1(_02727_),
    .A2(_02730_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15230_ (.A1(_02651_),
    .A2(\register_file[20][19] ),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15231_ (.I(_01083_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15232_ (.A1(_02403_),
    .A2(\register_file[21][19] ),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15233_ (.A1(_02732_),
    .A2(_02733_),
    .A3(_02734_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15234_ (.I(_01071_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15235_ (.A1(_02736_),
    .A2(\register_file[22][19] ),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15236_ (.I(_01325_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15237_ (.A1(_02488_),
    .A2(\register_file[23][19] ),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15238_ (.A1(_02737_),
    .A2(_02738_),
    .A3(_02739_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15239_ (.A1(_02735_),
    .A2(_02740_),
    .A3(_02658_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15240_ (.A1(_02731_),
    .A2(_02741_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15241_ (.A1(_02411_),
    .A2(\register_file[24][19] ),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15242_ (.A1(_02576_),
    .A2(\register_file[25][19] ),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15243_ (.A1(_02743_),
    .A2(_02744_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15244_ (.I(_01114_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15245_ (.A1(_02745_),
    .A2(_02746_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15246_ (.A1(_02747_),
    .A2(_01225_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15247_ (.A1(_02581_),
    .A2(\register_file[27][19] ),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15248_ (.A1(_02667_),
    .A2(\register_file[26][19] ),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15249_ (.I(_01075_),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15250_ (.A1(_02749_),
    .A2(_02750_),
    .B(_02751_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15251_ (.A1(_02748_),
    .A2(_02752_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15252_ (.A1(_02586_),
    .A2(\register_file[28][19] ),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15253_ (.A1(_02673_),
    .A2(\register_file[29][19] ),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15254_ (.A1(_02754_),
    .A2(_02672_),
    .A3(_02755_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15255_ (.A1(_02590_),
    .A2(\register_file[30][19] ),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15256_ (.A1(_02593_),
    .A2(\register_file[31][19] ),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15257_ (.A1(_02757_),
    .A2(_02592_),
    .A3(_02758_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15258_ (.A1(_02756_),
    .A2(_02759_),
    .A3(_02508_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15259_ (.A1(_02753_),
    .A2(_02760_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15260_ (.I(_01104_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15261_ (.A1(_02742_),
    .A2(_02761_),
    .A3(_02762_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15262_ (.I(_01079_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15263_ (.A1(_02764_),
    .A2(\register_file[8][19] ),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15264_ (.A1(_02513_),
    .A2(\register_file[9][19] ),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15265_ (.A1(_02765_),
    .A2(_02766_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15266_ (.A1(_02767_),
    .A2(_02685_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15267_ (.A1(_02768_),
    .A2(_02687_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15268_ (.A1(_02518_),
    .A2(\register_file[11][19] ),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15269_ (.A1(_02520_),
    .A2(\register_file[10][19] ),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15270_ (.A1(_02770_),
    .A2(_02771_),
    .B(_02691_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15271_ (.A1(_02769_),
    .A2(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15272_ (.A1(_02524_),
    .A2(\register_file[12][19] ),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15273_ (.A1(_02610_),
    .A2(\register_file[13][19] ),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15274_ (.A1(_02774_),
    .A2(_02609_),
    .A3(_02775_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15275_ (.A1(_02442_),
    .A2(\register_file[14][19] ),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15276_ (.A1(_02444_),
    .A2(\register_file[15][19] ),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15277_ (.A1(_02777_),
    .A2(_02529_),
    .A3(_02778_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15278_ (.A1(_02776_),
    .A2(_02779_),
    .A3(_02447_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15279_ (.A1(_02773_),
    .A2(_02780_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15280_ (.A1(_02450_),
    .A2(\register_file[6][19] ),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15281_ (.I(\register_file[7][19] ),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15282_ (.A1(_02783_),
    .A2(_02620_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15283_ (.A1(_02782_),
    .A2(_02784_),
    .A3(_02537_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15284_ (.I(_01530_),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15285_ (.I(\register_file[4][19] ),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15286_ (.A1(_02786_),
    .A2(_02787_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15287_ (.I(\register_file[5][19] ),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15288_ (.A1(_02789_),
    .A2(_02542_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15289_ (.A1(_02788_),
    .A2(_02790_),
    .A3(_02544_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15290_ (.A1(_02785_),
    .A2(_02791_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15291_ (.I(_01021_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15292_ (.A1(_02792_),
    .A2(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15293_ (.A1(_02548_),
    .A2(\register_file[2][19] ),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15294_ (.I(\register_file[3][19] ),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15295_ (.A1(_02796_),
    .A2(_02715_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15296_ (.A1(_02462_),
    .A2(_02795_),
    .A3(_02797_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15297_ (.A1(_02634_),
    .A2(\register_file[1][19] ),
    .B(_02635_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15298_ (.A1(_02798_),
    .A2(_02799_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15299_ (.I(_02800_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15300_ (.A1(_02794_),
    .A2(_02801_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15301_ (.A1(_02781_),
    .A2(_02802_),
    .A3(_02471_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15302_ (.A1(_02763_),
    .A2(_02803_),
    .B(_02473_),
    .ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15303_ (.A1(_02474_),
    .A2(\register_file[24][20] ),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15304_ (.I(_01058_),
    .Z(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15305_ (.A1(_02805_),
    .A2(\register_file[25][20] ),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15306_ (.A1(_02804_),
    .A2(_02806_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15307_ (.I(_01062_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15308_ (.A1(_02807_),
    .A2(_02808_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15309_ (.A1(_02809_),
    .A2(_01066_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15310_ (.A1(_02646_),
    .A2(\register_file[27][20] ),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15311_ (.I(_01042_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15312_ (.A1(_02812_),
    .A2(\register_file[26][20] ),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15313_ (.I(_01559_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15314_ (.A1(_02811_),
    .A2(_02813_),
    .B(_02814_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15315_ (.A1(_02810_),
    .A2(_02815_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15316_ (.A1(_02651_),
    .A2(\register_file[28][20] ),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15317_ (.I(_01038_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15318_ (.A1(_02818_),
    .A2(\register_file[29][20] ),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15319_ (.A1(_02817_),
    .A2(_02733_),
    .A3(_02819_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15320_ (.A1(_02736_),
    .A2(\register_file[30][20] ),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15321_ (.A1(_02488_),
    .A2(\register_file[31][20] ),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15322_ (.A1(_02821_),
    .A2(_02738_),
    .A3(_02822_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15323_ (.A1(_02820_),
    .A2(_02823_),
    .A3(_02658_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15324_ (.A1(_02816_),
    .A2(_02824_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15325_ (.I(_01107_),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15326_ (.A1(_02826_),
    .A2(\register_file[16][20] ),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15327_ (.A1(_02576_),
    .A2(\register_file[17][20] ),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15328_ (.A1(_02827_),
    .A2(_02828_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15329_ (.A1(_02829_),
    .A2(_02746_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15330_ (.A1(_02830_),
    .A2(_01010_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15331_ (.A1(_02581_),
    .A2(\register_file[19][20] ),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15332_ (.A1(_02667_),
    .A2(\register_file[18][20] ),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15333_ (.A1(_02832_),
    .A2(_02833_),
    .B(_02751_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15334_ (.A1(_02831_),
    .A2(_02834_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15335_ (.A1(_02586_),
    .A2(\register_file[20][20] ),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15336_ (.A1(_02673_),
    .A2(\register_file[21][20] ),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15337_ (.A1(_02836_),
    .A2(_02672_),
    .A3(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15338_ (.A1(_02590_),
    .A2(\register_file[22][20] ),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15339_ (.A1(_02593_),
    .A2(\register_file[23][20] ),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15340_ (.A1(_02839_),
    .A2(_02592_),
    .A3(_02840_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15341_ (.A1(_02838_),
    .A2(_02841_),
    .A3(_02508_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15342_ (.A1(_02835_),
    .A2(_02842_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15343_ (.A1(_02825_),
    .A2(_02843_),
    .A3(_02762_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15344_ (.A1(_02764_),
    .A2(\register_file[8][20] ),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15345_ (.A1(_02513_),
    .A2(\register_file[9][20] ),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15346_ (.A1(_02845_),
    .A2(_02846_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15347_ (.A1(_02847_),
    .A2(_02685_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15348_ (.A1(_02848_),
    .A2(_02687_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15349_ (.A1(_02518_),
    .A2(\register_file[11][20] ),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15350_ (.A1(_02520_),
    .A2(\register_file[10][20] ),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15351_ (.A1(_02850_),
    .A2(_02851_),
    .B(_02691_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15352_ (.A1(_02849_),
    .A2(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15353_ (.A1(_02524_),
    .A2(\register_file[12][20] ),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15354_ (.A1(_02610_),
    .A2(\register_file[13][20] ),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15355_ (.A1(_02854_),
    .A2(_02609_),
    .A3(_02855_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15356_ (.I(_01161_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15357_ (.A1(_02857_),
    .A2(\register_file[14][20] ),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15358_ (.I(_01455_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15359_ (.A1(_02859_),
    .A2(\register_file[15][20] ),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15360_ (.A1(_02858_),
    .A2(_02529_),
    .A3(_02860_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15361_ (.I(_01147_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15362_ (.A1(_02856_),
    .A2(_02861_),
    .A3(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15363_ (.A1(_02853_),
    .A2(_02863_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15364_ (.I(_01178_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15365_ (.A1(_02865_),
    .A2(\register_file[6][20] ),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15366_ (.I(\register_file[7][20] ),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15367_ (.A1(_02867_),
    .A2(_02620_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15368_ (.A1(_02866_),
    .A2(_02868_),
    .A3(_02537_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15369_ (.I(\register_file[4][20] ),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15370_ (.A1(_02786_),
    .A2(_02870_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15371_ (.I(\register_file[5][20] ),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15372_ (.A1(_02872_),
    .A2(_02542_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15373_ (.A1(_02871_),
    .A2(_02873_),
    .A3(_02544_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15374_ (.A1(_02869_),
    .A2(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15375_ (.A1(_02875_),
    .A2(_02793_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15376_ (.I(_01175_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15377_ (.A1(_02548_),
    .A2(\register_file[2][20] ),
    .Z(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15378_ (.I(\register_file[3][20] ),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15379_ (.A1(_02879_),
    .A2(_02715_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15380_ (.A1(_02877_),
    .A2(_02878_),
    .A3(_02880_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15381_ (.A1(_02634_),
    .A2(\register_file[1][20] ),
    .B(_02635_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15382_ (.A1(_02881_),
    .A2(_02882_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15383_ (.I(_02883_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15384_ (.A1(_02876_),
    .A2(_02884_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15385_ (.I(_01193_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15386_ (.A1(_02864_),
    .A2(_02885_),
    .A3(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15387_ (.I(_01199_),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15388_ (.A1(_02844_),
    .A2(_02887_),
    .B(_02888_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15389_ (.I(_01055_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15390_ (.A1(_02889_),
    .A2(\register_file[16][21] ),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15391_ (.A1(_02805_),
    .A2(\register_file[17][21] ),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15392_ (.A1(_02890_),
    .A2(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15393_ (.A1(_02892_),
    .A2(_02808_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15394_ (.A1(_02893_),
    .A2(_01292_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15395_ (.A1(_02646_),
    .A2(\register_file[19][21] ),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15396_ (.A1(_02812_),
    .A2(\register_file[18][21] ),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15397_ (.A1(_02895_),
    .A2(_02896_),
    .B(_02814_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15398_ (.A1(_02894_),
    .A2(_02897_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15399_ (.A1(_02651_),
    .A2(\register_file[20][21] ),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15400_ (.A1(_02818_),
    .A2(\register_file[21][21] ),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15401_ (.A1(_02899_),
    .A2(_02733_),
    .A3(_02900_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15402_ (.A1(_02736_),
    .A2(\register_file[22][21] ),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15403_ (.I(_01649_),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15404_ (.A1(_02903_),
    .A2(\register_file[23][21] ),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15405_ (.A1(_02902_),
    .A2(_02738_),
    .A3(_02904_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15406_ (.A1(_02901_),
    .A2(_02905_),
    .A3(_02658_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15407_ (.A1(_02898_),
    .A2(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15408_ (.A1(_02826_),
    .A2(\register_file[24][21] ),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15409_ (.A1(_02576_),
    .A2(\register_file[25][21] ),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15410_ (.A1(_02908_),
    .A2(_02909_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15411_ (.A1(_02910_),
    .A2(_02746_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15412_ (.I(_01065_),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15413_ (.A1(_02911_),
    .A2(_02912_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15414_ (.A1(_02581_),
    .A2(\register_file[27][21] ),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15415_ (.A1(_02667_),
    .A2(\register_file[26][21] ),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15416_ (.A1(_02914_),
    .A2(_02915_),
    .B(_02751_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15417_ (.A1(_02913_),
    .A2(_02916_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15418_ (.A1(_02586_),
    .A2(\register_file[28][21] ),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15419_ (.A1(_02673_),
    .A2(\register_file[29][21] ),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15420_ (.A1(_02918_),
    .A2(_02672_),
    .A3(_02919_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15421_ (.A1(_02590_),
    .A2(\register_file[30][21] ),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15422_ (.A1(_02593_),
    .A2(\register_file[31][21] ),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15423_ (.A1(_02921_),
    .A2(_02592_),
    .A3(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15424_ (.I(_01670_),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15425_ (.A1(_02920_),
    .A2(_02923_),
    .A3(_02924_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15426_ (.A1(_02917_),
    .A2(_02925_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15427_ (.A1(_02907_),
    .A2(_02926_),
    .A3(_02762_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15428_ (.A1(_02764_),
    .A2(\register_file[8][21] ),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15429_ (.I(_01013_),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15430_ (.A1(_02929_),
    .A2(\register_file[9][21] ),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15431_ (.A1(_02928_),
    .A2(_02930_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15432_ (.A1(_02931_),
    .A2(_02685_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15433_ (.A1(_02932_),
    .A2(_02687_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15434_ (.I(_01681_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15435_ (.A1(_02934_),
    .A2(\register_file[11][21] ),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15436_ (.I(_01138_),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15437_ (.A1(_02936_),
    .A2(\register_file[10][21] ),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15438_ (.A1(_02935_),
    .A2(_02937_),
    .B(_02691_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15439_ (.A1(_02933_),
    .A2(_02938_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15440_ (.I(_01018_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15441_ (.A1(_02940_),
    .A2(\register_file[12][21] ),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15442_ (.A1(_02610_),
    .A2(\register_file[13][21] ),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15443_ (.A1(_02941_),
    .A2(_02609_),
    .A3(_02942_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15444_ (.A1(_02857_),
    .A2(\register_file[14][21] ),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15445_ (.I(_01693_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15446_ (.A1(_02859_),
    .A2(\register_file[15][21] ),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15447_ (.A1(_02944_),
    .A2(_02945_),
    .A3(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15448_ (.A1(_02943_),
    .A2(_02947_),
    .A3(_02862_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15449_ (.A1(_02939_),
    .A2(_02948_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15450_ (.A1(_02865_),
    .A2(\register_file[6][21] ),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15451_ (.I(\register_file[7][21] ),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15452_ (.A1(_02951_),
    .A2(_02620_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15453_ (.I(_01092_),
    .Z(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15454_ (.A1(_02950_),
    .A2(_02952_),
    .A3(_02953_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15455_ (.I(\register_file[4][21] ),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15456_ (.A1(_02786_),
    .A2(_02955_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15457_ (.I(\register_file[5][21] ),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15458_ (.I(_00999_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15459_ (.A1(_02957_),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15460_ (.I(_01034_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15461_ (.A1(_02956_),
    .A2(_02959_),
    .A3(_02960_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15462_ (.A1(_02954_),
    .A2(_02961_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15463_ (.A1(_02962_),
    .A2(_02793_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15464_ (.I(_01151_),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15465_ (.A1(_02964_),
    .A2(\register_file[2][21] ),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15466_ (.I(\register_file[3][21] ),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15467_ (.A1(_02966_),
    .A2(_02715_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15468_ (.A1(_02877_),
    .A2(_02965_),
    .A3(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15469_ (.A1(_02634_),
    .A2(\register_file[1][21] ),
    .B(_02635_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15470_ (.A1(_02968_),
    .A2(_02969_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15471_ (.I(_02970_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15472_ (.A1(_02963_),
    .A2(_02971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15473_ (.A1(_02949_),
    .A2(_02972_),
    .A3(_02886_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15474_ (.A1(_02927_),
    .A2(_02973_),
    .B(_02888_),
    .ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15475_ (.A1(_02889_),
    .A2(\register_file[16][22] ),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15476_ (.A1(_02805_),
    .A2(\register_file[17][22] ),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15477_ (.A1(_02974_),
    .A2(_02975_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15478_ (.A1(_02976_),
    .A2(_02808_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15479_ (.I(_01009_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15480_ (.A1(_02977_),
    .A2(_02978_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15481_ (.A1(_02646_),
    .A2(\register_file[19][22] ),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15482_ (.A1(_02812_),
    .A2(\register_file[18][22] ),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15483_ (.A1(_02980_),
    .A2(_02981_),
    .B(_02814_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15484_ (.A1(_02979_),
    .A2(_02982_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15485_ (.A1(_02651_),
    .A2(\register_file[20][22] ),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15486_ (.A1(_02818_),
    .A2(\register_file[21][22] ),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15487_ (.A1(_02984_),
    .A2(_02733_),
    .A3(_02985_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15488_ (.A1(_02736_),
    .A2(\register_file[22][22] ),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15489_ (.A1(_02903_),
    .A2(\register_file[23][22] ),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15490_ (.A1(_02987_),
    .A2(_02738_),
    .A3(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15491_ (.A1(_02986_),
    .A2(_02989_),
    .A3(_02658_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15492_ (.A1(_02983_),
    .A2(_02990_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15493_ (.A1(_02826_),
    .A2(\register_file[24][22] ),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15494_ (.I(_01307_),
    .Z(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15495_ (.A1(_02993_),
    .A2(\register_file[25][22] ),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15496_ (.A1(_02992_),
    .A2(_02994_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15497_ (.A1(_02995_),
    .A2(_02746_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15498_ (.A1(_02996_),
    .A2(_02912_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15499_ (.I(_01119_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15500_ (.A1(_02998_),
    .A2(\register_file[27][22] ),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15501_ (.A1(_02667_),
    .A2(\register_file[26][22] ),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15502_ (.A1(_02999_),
    .A2(_03000_),
    .B(_02751_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15503_ (.A1(_02997_),
    .A2(_03001_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15504_ (.I(_01318_),
    .Z(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15505_ (.A1(_03003_),
    .A2(\register_file[28][22] ),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15506_ (.A1(_02673_),
    .A2(\register_file[29][22] ),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15507_ (.A1(_03004_),
    .A2(_02672_),
    .A3(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15508_ (.I(_01122_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15509_ (.A1(_03007_),
    .A2(\register_file[30][22] ),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15510_ (.I(_01093_),
    .Z(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15511_ (.I(_01142_),
    .Z(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15512_ (.A1(_03010_),
    .A2(\register_file[31][22] ),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15513_ (.A1(_03008_),
    .A2(_03009_),
    .A3(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15514_ (.A1(_03006_),
    .A2(_03012_),
    .A3(_02924_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15515_ (.A1(_03002_),
    .A2(_03013_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15516_ (.A1(_02991_),
    .A2(_03014_),
    .A3(_02762_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15517_ (.A1(_02764_),
    .A2(\register_file[8][22] ),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15518_ (.A1(_02929_),
    .A2(\register_file[9][22] ),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15519_ (.A1(_03016_),
    .A2(_03017_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15520_ (.A1(_03018_),
    .A2(_02685_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15521_ (.A1(_03019_),
    .A2(_02687_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15522_ (.A1(_02934_),
    .A2(\register_file[11][22] ),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15523_ (.A1(_02936_),
    .A2(\register_file[10][22] ),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15524_ (.A1(_03021_),
    .A2(_03022_),
    .B(_02691_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15525_ (.A1(_03020_),
    .A2(_03023_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15526_ (.A1(_02940_),
    .A2(\register_file[12][22] ),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15527_ (.I(_01774_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15528_ (.I(_01047_),
    .Z(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15529_ (.A1(_03027_),
    .A2(\register_file[13][22] ),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15530_ (.A1(_03025_),
    .A2(_03026_),
    .A3(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15531_ (.A1(_02857_),
    .A2(\register_file[14][22] ),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15532_ (.A1(_02859_),
    .A2(\register_file[15][22] ),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15533_ (.A1(_03030_),
    .A2(_02945_),
    .A3(_03031_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15534_ (.A1(_03029_),
    .A2(_03032_),
    .A3(_02862_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15535_ (.A1(_03024_),
    .A2(_03033_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15536_ (.A1(_02865_),
    .A2(\register_file[6][22] ),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15537_ (.I(\register_file[7][22] ),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15538_ (.I(_01354_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15539_ (.A1(_03036_),
    .A2(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15540_ (.A1(_03035_),
    .A2(_03038_),
    .A3(_02953_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15541_ (.I(\register_file[4][22] ),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15542_ (.A1(_02786_),
    .A2(_03040_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15543_ (.I(\register_file[5][22] ),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15544_ (.A1(_03042_),
    .A2(_02958_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15545_ (.A1(_03041_),
    .A2(_03043_),
    .A3(_02960_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15546_ (.A1(_03039_),
    .A2(_03044_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15547_ (.A1(_03045_),
    .A2(_02793_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15548_ (.A1(_02964_),
    .A2(\register_file[2][22] ),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15549_ (.I(\register_file[3][22] ),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15550_ (.A1(_03048_),
    .A2(_02715_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15551_ (.A1(_02877_),
    .A2(_03047_),
    .A3(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15552_ (.I(_01004_),
    .Z(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15553_ (.I(_01187_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15554_ (.A1(_03051_),
    .A2(\register_file[1][22] ),
    .B(_03052_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15555_ (.A1(_03050_),
    .A2(_03053_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15556_ (.I(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15557_ (.A1(_03046_),
    .A2(_03055_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15558_ (.A1(_03034_),
    .A2(_03056_),
    .A3(_02886_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15559_ (.A1(_03015_),
    .A2(_03057_),
    .B(_02888_),
    .ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15560_ (.A1(_02889_),
    .A2(\register_file[24][23] ),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15561_ (.A1(_02805_),
    .A2(\register_file[25][23] ),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15562_ (.A1(_03058_),
    .A2(_03059_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15563_ (.A1(_03060_),
    .A2(_02808_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15564_ (.A1(_03061_),
    .A2(_01066_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15565_ (.I(_01068_),
    .Z(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15566_ (.A1(_03063_),
    .A2(\register_file[27][23] ),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15567_ (.A1(_02812_),
    .A2(\register_file[26][23] ),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15568_ (.A1(_03064_),
    .A2(_03065_),
    .B(_02814_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15569_ (.A1(_03062_),
    .A2(_03066_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15570_ (.I(_01080_),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15571_ (.A1(_03068_),
    .A2(\register_file[28][23] ),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15572_ (.A1(_02818_),
    .A2(\register_file[29][23] ),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15573_ (.A1(_03069_),
    .A2(_02733_),
    .A3(_03070_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15574_ (.A1(_02736_),
    .A2(\register_file[30][23] ),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15575_ (.A1(_02903_),
    .A2(\register_file[31][23] ),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15576_ (.A1(_03072_),
    .A2(_02738_),
    .A3(_03073_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15577_ (.I(_01100_),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15578_ (.A1(_03071_),
    .A2(_03074_),
    .A3(_03075_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15579_ (.A1(_03067_),
    .A2(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15580_ (.A1(_02826_),
    .A2(\register_file[16][23] ),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15581_ (.A1(_02993_),
    .A2(\register_file[17][23] ),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15582_ (.A1(_03078_),
    .A2(_03079_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15583_ (.A1(_03080_),
    .A2(_02746_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15584_ (.A1(_03081_),
    .A2(_01010_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15585_ (.A1(_02998_),
    .A2(\register_file[19][23] ),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15586_ (.I(_01404_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15587_ (.A1(_03084_),
    .A2(\register_file[18][23] ),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15588_ (.A1(_03083_),
    .A2(_03085_),
    .B(_02751_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15589_ (.A1(_03082_),
    .A2(_03086_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15590_ (.A1(_03003_),
    .A2(\register_file[20][23] ),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15591_ (.I(_01132_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15592_ (.I(_01134_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15593_ (.A1(_03090_),
    .A2(\register_file[21][23] ),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15594_ (.A1(_03088_),
    .A2(_03089_),
    .A3(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15595_ (.A1(_03007_),
    .A2(\register_file[22][23] ),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15596_ (.A1(_03010_),
    .A2(\register_file[23][23] ),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15597_ (.A1(_03093_),
    .A2(_03009_),
    .A3(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15598_ (.A1(_03092_),
    .A2(_03095_),
    .A3(_02924_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15599_ (.A1(_03087_),
    .A2(_03096_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15600_ (.A1(_03077_),
    .A2(_03097_),
    .A3(_02762_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15601_ (.A1(_02764_),
    .A2(\register_file[8][23] ),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15602_ (.A1(_02929_),
    .A2(\register_file[9][23] ),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15603_ (.A1(_03099_),
    .A2(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15604_ (.I(_01423_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15605_ (.A1(_03101_),
    .A2(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15606_ (.I(_01426_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15607_ (.A1(_03103_),
    .A2(_03104_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15608_ (.A1(_02934_),
    .A2(\register_file[11][23] ),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15609_ (.A1(_02936_),
    .A2(\register_file[10][23] ),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15610_ (.I(_01074_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15611_ (.A1(_03106_),
    .A2(_03107_),
    .B(_03108_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15612_ (.D(_00000_),
    .CLK(clknet_leaf_37_clk),
    .Q(\register_file[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15613_ (.D(_00001_),
    .CLK(clknet_leaf_32_clk),
    .Q(\register_file[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15614_ (.D(_00002_),
    .CLK(clknet_leaf_24_clk),
    .Q(\register_file[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15615_ (.D(_00003_),
    .CLK(clknet_leaf_19_clk),
    .Q(\register_file[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15616_ (.D(_00004_),
    .CLK(clknet_leaf_19_clk),
    .Q(\register_file[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15617_ (.D(_00005_),
    .CLK(clknet_leaf_19_clk),
    .Q(\register_file[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15618_ (.D(_00006_),
    .CLK(clknet_leaf_20_clk),
    .Q(\register_file[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15619_ (.D(_00007_),
    .CLK(clknet_leaf_20_clk),
    .Q(\register_file[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15620_ (.D(_00008_),
    .CLK(clknet_leaf_72_clk),
    .Q(\register_file[30][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15621_ (.D(_00009_),
    .CLK(clknet_leaf_72_clk),
    .Q(\register_file[30][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15622_ (.D(_00010_),
    .CLK(clknet_leaf_89_clk),
    .Q(\register_file[30][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15623_ (.D(_00011_),
    .CLK(clknet_leaf_88_clk),
    .Q(\register_file[30][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15624_ (.D(_00012_),
    .CLK(clknet_leaf_89_clk),
    .Q(\register_file[30][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15625_ (.D(_00013_),
    .CLK(clknet_leaf_100_clk),
    .Q(\register_file[30][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15626_ (.D(_00014_),
    .CLK(clknet_leaf_99_clk),
    .Q(\register_file[30][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15627_ (.D(_00015_),
    .CLK(clknet_leaf_99_clk),
    .Q(\register_file[30][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15628_ (.D(_00016_),
    .CLK(clknet_leaf_135_clk),
    .Q(\register_file[30][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15629_ (.D(_00017_),
    .CLK(clknet_leaf_135_clk),
    .Q(\register_file[30][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15630_ (.D(_00018_),
    .CLK(clknet_leaf_152_clk),
    .Q(\register_file[30][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15631_ (.D(_00019_),
    .CLK(clknet_leaf_152_clk),
    .Q(\register_file[30][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15632_ (.D(_00020_),
    .CLK(clknet_leaf_165_clk),
    .Q(\register_file[30][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15633_ (.D(_00021_),
    .CLK(clknet_leaf_165_clk),
    .Q(\register_file[30][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15634_ (.D(_00022_),
    .CLK(clknet_leaf_178_clk),
    .Q(\register_file[30][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15635_ (.D(_00023_),
    .CLK(clknet_leaf_178_clk),
    .Q(\register_file[30][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15636_ (.D(_00024_),
    .CLK(clknet_leaf_210_clk),
    .Q(\register_file[30][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15637_ (.D(_00025_),
    .CLK(clknet_leaf_211_clk),
    .Q(\register_file[30][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15638_ (.D(_00026_),
    .CLK(clknet_leaf_212_clk),
    .Q(\register_file[30][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15639_ (.D(_00027_),
    .CLK(clknet_leaf_212_clk),
    .Q(\register_file[30][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15640_ (.D(_00028_),
    .CLK(clknet_leaf_197_clk),
    .Q(\register_file[30][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15641_ (.D(_00029_),
    .CLK(clknet_leaf_199_clk),
    .Q(\register_file[30][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15642_ (.D(_00030_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\register_file[30][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15643_ (.D(_00031_),
    .CLK(clknet_leaf_271_clk),
    .Q(\register_file[30][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15644_ (.D(_00032_),
    .CLK(clknet_leaf_282_clk),
    .Q(\register_file[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15645_ (.D(_00033_),
    .CLK(clknet_leaf_302_clk),
    .Q(\register_file[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15646_ (.D(_00034_),
    .CLK(clknet_leaf_304_clk),
    .Q(\register_file[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15647_ (.D(_00035_),
    .CLK(clknet_leaf_3_clk),
    .Q(\register_file[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15648_ (.D(_00036_),
    .CLK(clknet_leaf_3_clk),
    .Q(\register_file[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15649_ (.D(_00037_),
    .CLK(clknet_leaf_20_clk),
    .Q(\register_file[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15650_ (.D(_00038_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\register_file[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15651_ (.D(_00039_),
    .CLK(clknet_leaf_53_clk),
    .Q(\register_file[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15652_ (.D(_00040_),
    .CLK(clknet_leaf_69_clk),
    .Q(\register_file[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15653_ (.D(_00041_),
    .CLK(clknet_leaf_69_clk),
    .Q(\register_file[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15654_ (.D(_00042_),
    .CLK(clknet_leaf_88_clk),
    .Q(\register_file[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15655_ (.D(_00043_),
    .CLK(clknet_leaf_88_clk),
    .Q(\register_file[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15656_ (.D(_00044_),
    .CLK(clknet_leaf_94_clk),
    .Q(\register_file[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15657_ (.D(_00045_),
    .CLK(clknet_leaf_94_clk),
    .Q(\register_file[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15658_ (.D(_00046_),
    .CLK(clknet_leaf_94_clk),
    .Q(\register_file[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15659_ (.D(_00047_),
    .CLK(clknet_leaf_141_clk),
    .Q(\register_file[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15660_ (.D(_00048_),
    .CLK(clknet_leaf_135_clk),
    .Q(\register_file[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15661_ (.D(_00049_),
    .CLK(clknet_leaf_142_clk),
    .Q(\register_file[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15662_ (.D(_00050_),
    .CLK(clknet_leaf_147_clk),
    .Q(\register_file[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15663_ (.D(_00051_),
    .CLK(clknet_leaf_146_clk),
    .Q(\register_file[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15664_ (.D(_00052_),
    .CLK(clknet_leaf_173_clk),
    .Q(\register_file[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15665_ (.D(_00053_),
    .CLK(clknet_leaf_173_clk),
    .Q(\register_file[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15666_ (.D(_00054_),
    .CLK(clknet_leaf_178_clk),
    .Q(\register_file[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15667_ (.D(_00055_),
    .CLK(clknet_leaf_210_clk),
    .Q(\register_file[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15668_ (.D(_00056_),
    .CLK(clknet_leaf_210_clk),
    .Q(\register_file[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15669_ (.D(_00057_),
    .CLK(clknet_leaf_224_clk),
    .Q(\register_file[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15670_ (.D(_00058_),
    .CLK(clknet_leaf_225_clk),
    .Q(\register_file[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15671_ (.D(_00059_),
    .CLK(clknet_leaf_224_clk),
    .Q(\register_file[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15672_ (.D(_00060_),
    .CLK(clknet_leaf_240_clk),
    .Q(\register_file[2][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15673_ (.D(_00061_),
    .CLK(clknet_leaf_241_clk),
    .Q(\register_file[2][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15674_ (.D(_00062_),
    .CLK(clknet_leaf_257_clk),
    .Q(\register_file[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15675_ (.D(_00063_),
    .CLK(clknet_leaf_284_clk),
    .Q(\register_file[2][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15676_ (.D(_00064_),
    .CLK(clknet_leaf_36_clk),
    .Q(\register_file[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15677_ (.D(_00065_),
    .CLK(clknet_leaf_32_clk),
    .Q(\register_file[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15678_ (.D(_00066_),
    .CLK(clknet_leaf_24_clk),
    .Q(\register_file[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15679_ (.D(_00067_),
    .CLK(clknet_leaf_19_clk),
    .Q(\register_file[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15680_ (.D(_00068_),
    .CLK(clknet_leaf_16_clk),
    .Q(\register_file[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15681_ (.D(_00069_),
    .CLK(clknet_leaf_19_clk),
    .Q(\register_file[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15682_ (.D(_00070_),
    .CLK(clknet_leaf_19_clk),
    .Q(\register_file[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15683_ (.D(_00071_),
    .CLK(clknet_leaf_20_clk),
    .Q(\register_file[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15684_ (.D(_00072_),
    .CLK(clknet_leaf_70_clk),
    .Q(\register_file[28][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15685_ (.D(_00073_),
    .CLK(clknet_leaf_72_clk),
    .Q(\register_file[28][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15686_ (.D(_00074_),
    .CLK(clknet_leaf_83_clk),
    .Q(\register_file[28][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15687_ (.D(_00075_),
    .CLK(clknet_leaf_85_clk),
    .Q(\register_file[28][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15688_ (.D(_00076_),
    .CLK(clknet_leaf_84_clk),
    .Q(\register_file[28][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15689_ (.D(_00077_),
    .CLK(clknet_leaf_101_clk),
    .Q(\register_file[28][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15690_ (.D(_00078_),
    .CLK(clknet_leaf_100_clk),
    .Q(\register_file[28][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15691_ (.D(_00079_),
    .CLK(clknet_leaf_135_clk),
    .Q(\register_file[28][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15692_ (.D(_00080_),
    .CLK(clknet_leaf_134_clk),
    .Q(\register_file[28][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15693_ (.D(_00081_),
    .CLK(clknet_leaf_148_clk),
    .Q(\register_file[28][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15694_ (.D(_00082_),
    .CLK(clknet_leaf_152_clk),
    .Q(\register_file[28][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15695_ (.D(_00083_),
    .CLK(clknet_leaf_152_clk),
    .Q(\register_file[28][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15696_ (.D(_00084_),
    .CLK(clknet_leaf_165_clk),
    .Q(\register_file[28][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15697_ (.D(_00085_),
    .CLK(clknet_leaf_166_clk),
    .Q(\register_file[28][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15698_ (.D(_00086_),
    .CLK(clknet_leaf_178_clk),
    .Q(\register_file[28][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15699_ (.D(_00087_),
    .CLK(clknet_leaf_179_clk),
    .Q(\register_file[28][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15700_ (.D(_00088_),
    .CLK(clknet_leaf_179_clk),
    .Q(\register_file[28][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15701_ (.D(_00089_),
    .CLK(clknet_leaf_211_clk),
    .Q(\register_file[28][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15702_ (.D(_00090_),
    .CLK(clknet_leaf_212_clk),
    .Q(\register_file[28][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15703_ (.D(_00091_),
    .CLK(clknet_leaf_212_clk),
    .Q(\register_file[28][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15704_ (.D(_00092_),
    .CLK(clknet_leaf_196_clk),
    .Q(\register_file[28][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15705_ (.D(_00093_),
    .CLK(clknet_leaf_199_clk),
    .Q(\register_file[28][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15706_ (.D(_00094_),
    .CLK(clknet_leaf_267_clk),
    .Q(\register_file[28][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15707_ (.D(_00095_),
    .CLK(clknet_leaf_271_clk),
    .Q(\register_file[28][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15708_ (.D(_00096_),
    .CLK(clknet_leaf_36_clk),
    .Q(\register_file[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15709_ (.D(_00097_),
    .CLK(clknet_leaf_32_clk),
    .Q(\register_file[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15710_ (.D(_00098_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\register_file[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15711_ (.D(_00099_),
    .CLK(clknet_leaf_15_clk),
    .Q(\register_file[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15712_ (.D(_00100_),
    .CLK(clknet_leaf_15_clk),
    .Q(\register_file[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15713_ (.D(_00101_),
    .CLK(clknet_leaf_53_clk),
    .Q(\register_file[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15714_ (.D(_00102_),
    .CLK(clknet_leaf_54_clk),
    .Q(\register_file[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15715_ (.D(_00103_),
    .CLK(clknet_leaf_54_clk),
    .Q(\register_file[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15716_ (.D(_00104_),
    .CLK(clknet_leaf_70_clk),
    .Q(\register_file[27][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15717_ (.D(_00105_),
    .CLK(clknet_leaf_69_clk),
    .Q(\register_file[27][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15718_ (.D(_00106_),
    .CLK(clknet_leaf_88_clk),
    .Q(\register_file[27][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15719_ (.D(_00107_),
    .CLK(clknet_leaf_88_clk),
    .Q(\register_file[27][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15720_ (.D(_00108_),
    .CLK(clknet_leaf_88_clk),
    .Q(\register_file[27][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15721_ (.D(_00109_),
    .CLK(clknet_leaf_94_clk),
    .Q(\register_file[27][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15722_ (.D(_00110_),
    .CLK(clknet_leaf_101_clk),
    .Q(\register_file[27][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15723_ (.D(_00111_),
    .CLK(clknet_leaf_136_clk),
    .Q(\register_file[27][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15724_ (.D(_00112_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\register_file[27][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15725_ (.D(_00113_),
    .CLK(clknet_leaf_136_clk),
    .Q(\register_file[27][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15726_ (.D(_00114_),
    .CLK(clknet_leaf_146_clk),
    .Q(\register_file[27][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15727_ (.D(_00115_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\register_file[27][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15728_ (.D(_00116_),
    .CLK(clknet_leaf_166_clk),
    .Q(\register_file[27][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15729_ (.D(_00117_),
    .CLK(clknet_leaf_166_clk),
    .Q(\register_file[27][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15730_ (.D(_00118_),
    .CLK(clknet_leaf_173_clk),
    .Q(\register_file[27][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15731_ (.D(_00119_),
    .CLK(clknet_leaf_177_clk),
    .Q(\register_file[27][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15732_ (.D(_00120_),
    .CLK(clknet_leaf_177_clk),
    .Q(\register_file[27][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15733_ (.D(_00121_),
    .CLK(clknet_leaf_211_clk),
    .Q(\register_file[27][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15734_ (.D(_00122_),
    .CLK(clknet_leaf_212_clk),
    .Q(\register_file[27][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15735_ (.D(_00123_),
    .CLK(clknet_leaf_212_clk),
    .Q(\register_file[27][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15736_ (.D(_00124_),
    .CLK(clknet_leaf_199_clk),
    .Q(\register_file[27][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15737_ (.D(_00125_),
    .CLK(clknet_leaf_262_clk),
    .Q(\register_file[27][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15738_ (.D(_00126_),
    .CLK(clknet_leaf_267_clk),
    .Q(\register_file[27][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15739_ (.D(_00127_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\register_file[27][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15740_ (.D(_00128_),
    .CLK(clknet_leaf_283_clk),
    .Q(\register_file[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15741_ (.D(_00129_),
    .CLK(clknet_leaf_281_clk),
    .Q(\register_file[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15742_ (.D(_00130_),
    .CLK(clknet_leaf_8_clk),
    .Q(\register_file[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15743_ (.D(_00131_),
    .CLK(clknet_leaf_4_clk),
    .Q(\register_file[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15744_ (.D(_00132_),
    .CLK(clknet_leaf_4_clk),
    .Q(\register_file[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15745_ (.D(_00133_),
    .CLK(clknet_leaf_53_clk),
    .Q(\register_file[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15746_ (.D(_00134_),
    .CLK(clknet_leaf_53_clk),
    .Q(\register_file[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15747_ (.D(_00135_),
    .CLK(clknet_leaf_54_clk),
    .Q(\register_file[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15748_ (.D(_00136_),
    .CLK(clknet_leaf_69_clk),
    .Q(\register_file[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15749_ (.D(_00137_),
    .CLK(clknet_leaf_69_clk),
    .Q(\register_file[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15750_ (.D(_00138_),
    .CLK(clknet_leaf_83_clk),
    .Q(\register_file[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15751_ (.D(_00139_),
    .CLK(clknet_leaf_84_clk),
    .Q(\register_file[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15752_ (.D(_00140_),
    .CLK(clknet_leaf_84_clk),
    .Q(\register_file[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15753_ (.D(_00141_),
    .CLK(clknet_leaf_100_clk),
    .Q(\register_file[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15754_ (.D(_00142_),
    .CLK(clknet_leaf_95_clk),
    .Q(\register_file[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15755_ (.D(_00143_),
    .CLK(clknet_leaf_136_clk),
    .Q(\register_file[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15756_ (.D(_00144_),
    .CLK(clknet_leaf_136_clk),
    .Q(\register_file[13][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15757_ (.D(_00145_),
    .CLK(clknet_leaf_148_clk),
    .Q(\register_file[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15758_ (.D(_00146_),
    .CLK(clknet_leaf_148_clk),
    .Q(\register_file[13][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15759_ (.D(_00147_),
    .CLK(clknet_leaf_146_clk),
    .Q(\register_file[13][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15760_ (.D(_00148_),
    .CLK(clknet_leaf_173_clk),
    .Q(\register_file[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15761_ (.D(_00149_),
    .CLK(clknet_leaf_173_clk),
    .Q(\register_file[13][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15762_ (.D(_00150_),
    .CLK(clknet_leaf_177_clk),
    .Q(\register_file[13][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15763_ (.D(_00151_),
    .CLK(clknet_leaf_177_clk),
    .Q(\register_file[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15764_ (.D(_00152_),
    .CLK(clknet_leaf_177_clk),
    .Q(\register_file[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15765_ (.D(_00153_),
    .CLK(clknet_leaf_217_clk),
    .Q(\register_file[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15766_ (.D(_00154_),
    .CLK(clknet_leaf_224_clk),
    .Q(\register_file[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15767_ (.D(_00155_),
    .CLK(clknet_leaf_224_clk),
    .Q(\register_file[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15768_ (.D(_00156_),
    .CLK(clknet_leaf_259_clk),
    .Q(\register_file[13][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15769_ (.D(_00157_),
    .CLK(clknet_leaf_259_clk),
    .Q(\register_file[13][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15770_ (.D(_00158_),
    .CLK(clknet_leaf_255_clk),
    .Q(\register_file[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15771_ (.D(_00159_),
    .CLK(clknet_leaf_283_clk),
    .Q(\register_file[13][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15772_ (.D(_00160_),
    .CLK(clknet_leaf_279_clk),
    .Q(\register_file[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15773_ (.D(_00161_),
    .CLK(clknet_leaf_280_clk),
    .Q(\register_file[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15774_ (.D(_00162_),
    .CLK(clknet_leaf_29_clk),
    .Q(\register_file[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15775_ (.D(_00163_),
    .CLK(clknet_leaf_12_clk),
    .Q(\register_file[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15776_ (.D(_00164_),
    .CLK(clknet_leaf_13_clk),
    .Q(\register_file[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15777_ (.D(_00165_),
    .CLK(clknet_leaf_52_clk),
    .Q(\register_file[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15778_ (.D(_00166_),
    .CLK(clknet_leaf_52_clk),
    .Q(\register_file[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15779_ (.D(_00167_),
    .CLK(clknet_leaf_56_clk),
    .Q(\register_file[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15780_ (.D(_00168_),
    .CLK(clknet_leaf_66_clk),
    .Q(\register_file[19][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15781_ (.D(_00169_),
    .CLK(clknet_leaf_66_clk),
    .Q(\register_file[19][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15782_ (.D(_00170_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\register_file[19][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15783_ (.D(_00171_),
    .CLK(clknet_leaf_47_clk),
    .Q(\register_file[19][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15784_ (.D(_00172_),
    .CLK(clknet_leaf_108_clk),
    .Q(\register_file[19][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15785_ (.D(_00173_),
    .CLK(clknet_leaf_103_clk),
    .Q(\register_file[19][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15786_ (.D(_00174_),
    .CLK(clknet_leaf_103_clk),
    .Q(\register_file[19][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15787_ (.D(_00175_),
    .CLK(clknet_leaf_131_clk),
    .Q(\register_file[19][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15788_ (.D(_00176_),
    .CLK(clknet_leaf_123_clk),
    .Q(\register_file[19][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15789_ (.D(_00177_),
    .CLK(clknet_leaf_123_clk),
    .Q(\register_file[19][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15790_ (.D(_00178_),
    .CLK(clknet_leaf_127_clk),
    .Q(\register_file[19][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15791_ (.D(_00179_),
    .CLK(clknet_leaf_127_clk),
    .Q(\register_file[19][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15792_ (.D(_00180_),
    .CLK(clknet_leaf_169_clk),
    .Q(\register_file[19][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15793_ (.D(_00181_),
    .CLK(clknet_leaf_168_clk),
    .Q(\register_file[19][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15794_ (.D(_00182_),
    .CLK(clknet_leaf_168_clk),
    .Q(\register_file[19][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15795_ (.D(_00183_),
    .CLK(clknet_leaf_172_clk),
    .Q(\register_file[19][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15796_ (.D(_00184_),
    .CLK(clknet_leaf_172_clk),
    .Q(\register_file[19][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15797_ (.D(_00185_),
    .CLK(clknet_leaf_205_clk),
    .Q(\register_file[19][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15798_ (.D(_00186_),
    .CLK(clknet_leaf_204_clk),
    .Q(\register_file[19][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15799_ (.D(_00187_),
    .CLK(clknet_leaf_214_clk),
    .Q(\register_file[19][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15800_ (.D(_00188_),
    .CLK(clknet_leaf_261_clk),
    .Q(\register_file[19][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15801_ (.D(_00189_),
    .CLK(clknet_leaf_261_clk),
    .Q(\register_file[19][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15802_ (.D(_00190_),
    .CLK(clknet_leaf_276_clk),
    .Q(\register_file[19][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15803_ (.D(_00191_),
    .CLK(clknet_leaf_275_clk),
    .Q(\register_file[19][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15804_ (.D(_00192_),
    .CLK(clknet_leaf_276_clk),
    .Q(\register_file[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15805_ (.D(_00193_),
    .CLK(clknet_leaf_279_clk),
    .Q(\register_file[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15806_ (.D(_00194_),
    .CLK(clknet_leaf_28_clk),
    .Q(\register_file[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15807_ (.D(_00195_),
    .CLK(clknet_leaf_11_clk),
    .Q(\register_file[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15808_ (.D(_00196_),
    .CLK(clknet_leaf_10_clk),
    .Q(\register_file[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15809_ (.D(_00197_),
    .CLK(clknet_leaf_50_clk),
    .Q(\register_file[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15810_ (.D(_00198_),
    .CLK(clknet_leaf_49_clk),
    .Q(\register_file[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15811_ (.D(_00199_),
    .CLK(clknet_leaf_49_clk),
    .Q(\register_file[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15812_ (.D(_00200_),
    .CLK(clknet_leaf_62_clk),
    .Q(\register_file[26][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15813_ (.D(_00201_),
    .CLK(clknet_leaf_64_clk),
    .Q(\register_file[26][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15814_ (.D(_00202_),
    .CLK(clknet_leaf_107_clk),
    .Q(\register_file[26][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15815_ (.D(_00203_),
    .CLK(clknet_leaf_107_clk),
    .Q(\register_file[26][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15816_ (.D(_00204_),
    .CLK(clknet_leaf_107_clk),
    .Q(\register_file[26][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15817_ (.D(_00205_),
    .CLK(clknet_leaf_105_clk),
    .Q(\register_file[26][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15818_ (.D(_00206_),
    .CLK(clknet_leaf_104_clk),
    .Q(\register_file[26][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15819_ (.D(_00207_),
    .CLK(clknet_leaf_132_clk),
    .Q(\register_file[26][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15820_ (.D(_00208_),
    .CLK(clknet_leaf_132_clk),
    .Q(\register_file[26][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15821_ (.D(_00209_),
    .CLK(clknet_leaf_131_clk),
    .Q(\register_file[26][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15822_ (.D(_00210_),
    .CLK(clknet_leaf_150_clk),
    .Q(\register_file[26][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15823_ (.D(_00211_),
    .CLK(clknet_leaf_127_clk),
    .Q(\register_file[26][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15824_ (.D(_00212_),
    .CLK(clknet_leaf_169_clk),
    .Q(\register_file[26][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15825_ (.D(_00213_),
    .CLK(clknet_leaf_170_clk),
    .Q(\register_file[26][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15826_ (.D(_00214_),
    .CLK(clknet_leaf_169_clk),
    .Q(\register_file[26][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15827_ (.D(_00215_),
    .CLK(clknet_leaf_173_clk),
    .Q(\register_file[26][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15828_ (.D(_00216_),
    .CLK(clknet_leaf_172_clk),
    .Q(\register_file[26][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15829_ (.D(_00217_),
    .CLK(clknet_leaf_219_clk),
    .Q(\register_file[26][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15830_ (.D(_00218_),
    .CLK(clknet_leaf_219_clk),
    .Q(\register_file[26][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15831_ (.D(_00219_),
    .CLK(clknet_leaf_219_clk),
    .Q(\register_file[26][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15832_ (.D(_00220_),
    .CLK(clknet_leaf_260_clk),
    .Q(\register_file[26][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15833_ (.D(_00221_),
    .CLK(clknet_leaf_263_clk),
    .Q(\register_file[26][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15834_ (.D(_00222_),
    .CLK(clknet_leaf_265_clk),
    .Q(\register_file[26][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15835_ (.D(_00223_),
    .CLK(clknet_leaf_274_clk),
    .Q(\register_file[26][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15836_ (.D(_00224_),
    .CLK(clknet_leaf_279_clk),
    .Q(\register_file[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15837_ (.D(_00225_),
    .CLK(clknet_leaf_279_clk),
    .Q(\register_file[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15838_ (.D(_00226_),
    .CLK(clknet_leaf_8_clk),
    .Q(\register_file[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15839_ (.D(_00227_),
    .CLK(clknet_leaf_13_clk),
    .Q(\register_file[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15840_ (.D(_00228_),
    .CLK(clknet_leaf_5_clk),
    .Q(\register_file[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15841_ (.D(_00229_),
    .CLK(clknet_leaf_22_clk),
    .Q(\register_file[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15842_ (.D(_00230_),
    .CLK(clknet_leaf_52_clk),
    .Q(\register_file[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15843_ (.D(_00231_),
    .CLK(clknet_leaf_56_clk),
    .Q(\register_file[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15844_ (.D(_00232_),
    .CLK(clknet_leaf_61_clk),
    .Q(\register_file[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15845_ (.D(_00233_),
    .CLK(clknet_leaf_61_clk),
    .Q(\register_file[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15846_ (.D(_00234_),
    .CLK(clknet_leaf_47_clk),
    .Q(\register_file[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15847_ (.D(_00235_),
    .CLK(clknet_leaf_46_clk),
    .Q(\register_file[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15848_ (.D(_00236_),
    .CLK(clknet_leaf_108_clk),
    .Q(\register_file[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15849_ (.D(_00237_),
    .CLK(clknet_leaf_111_clk),
    .Q(\register_file[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15850_ (.D(_00238_),
    .CLK(clknet_leaf_111_clk),
    .Q(\register_file[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15851_ (.D(_00239_),
    .CLK(clknet_leaf_122_clk),
    .Q(\register_file[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15852_ (.D(_00240_),
    .CLK(clknet_leaf_122_clk),
    .Q(\register_file[12][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15853_ (.D(_00241_),
    .CLK(clknet_leaf_126_clk),
    .Q(\register_file[12][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15854_ (.D(_00242_),
    .CLK(clknet_leaf_126_clk),
    .Q(\register_file[12][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15855_ (.D(_00243_),
    .CLK(clknet_leaf_127_clk),
    .Q(\register_file[12][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15856_ (.D(_00244_),
    .CLK(clknet_leaf_170_clk),
    .Q(\register_file[12][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15857_ (.D(_00245_),
    .CLK(clknet_leaf_171_clk),
    .Q(\register_file[12][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15858_ (.D(_00246_),
    .CLK(clknet_leaf_171_clk),
    .Q(\register_file[12][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15859_ (.D(_00247_),
    .CLK(clknet_leaf_176_clk),
    .Q(\register_file[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15860_ (.D(_00248_),
    .CLK(clknet_leaf_175_clk),
    .Q(\register_file[12][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15861_ (.D(_00249_),
    .CLK(clknet_leaf_218_clk),
    .Q(\register_file[12][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15862_ (.D(_00250_),
    .CLK(clknet_leaf_220_clk),
    .Q(\register_file[12][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15863_ (.D(_00251_),
    .CLK(clknet_leaf_223_clk),
    .Q(\register_file[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15864_ (.D(_00252_),
    .CLK(clknet_leaf_260_clk),
    .Q(\register_file[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15865_ (.D(_00253_),
    .CLK(clknet_leaf_260_clk),
    .Q(\register_file[12][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15866_ (.D(_00254_),
    .CLK(clknet_leaf_255_clk),
    .Q(\register_file[12][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15867_ (.D(_00255_),
    .CLK(clknet_leaf_275_clk),
    .Q(\register_file[12][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15868_ (.D(_00256_),
    .CLK(clknet_leaf_276_clk),
    .Q(\register_file[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15869_ (.D(_00257_),
    .CLK(clknet_leaf_280_clk),
    .Q(\register_file[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15870_ (.D(_00258_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\register_file[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15871_ (.D(_00259_),
    .CLK(clknet_leaf_10_clk),
    .Q(\register_file[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15872_ (.D(_00260_),
    .CLK(clknet_leaf_7_clk),
    .Q(\register_file[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15873_ (.D(_00261_),
    .CLK(clknet_leaf_23_clk),
    .Q(\register_file[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15874_ (.D(_00262_),
    .CLK(clknet_leaf_50_clk),
    .Q(\register_file[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15875_ (.D(_00263_),
    .CLK(clknet_leaf_50_clk),
    .Q(\register_file[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15876_ (.D(_00264_),
    .CLK(clknet_leaf_62_clk),
    .Q(\register_file[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15877_ (.D(_00265_),
    .CLK(clknet_leaf_63_clk),
    .Q(\register_file[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15878_ (.D(_00266_),
    .CLK(clknet_leaf_46_clk),
    .Q(\register_file[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15879_ (.D(_00267_),
    .CLK(clknet_leaf_109_clk),
    .Q(\register_file[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15880_ (.D(_00268_),
    .CLK(clknet_leaf_109_clk),
    .Q(\register_file[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15881_ (.D(_00269_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\register_file[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15882_ (.D(_00270_),
    .CLK(clknet_leaf_112_clk),
    .Q(\register_file[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15883_ (.D(_00271_),
    .CLK(clknet_leaf_121_clk),
    .Q(\register_file[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15884_ (.D(_00272_),
    .CLK(clknet_leaf_124_clk),
    .Q(\register_file[11][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15885_ (.D(_00273_),
    .CLK(clknet_leaf_121_clk),
    .Q(\register_file[11][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15886_ (.D(_00274_),
    .CLK(clknet_leaf_187_clk),
    .Q(\register_file[11][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15887_ (.D(_00275_),
    .CLK(clknet_leaf_186_clk),
    .Q(\register_file[11][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15888_ (.D(_00276_),
    .CLK(clknet_leaf_186_clk),
    .Q(\register_file[11][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15889_ (.D(_00277_),
    .CLK(clknet_leaf_171_clk),
    .Q(\register_file[11][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15890_ (.D(_00278_),
    .CLK(clknet_leaf_171_clk),
    .Q(\register_file[11][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15891_ (.D(_00279_),
    .CLK(clknet_leaf_213_clk),
    .Q(\register_file[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15892_ (.D(_00280_),
    .CLK(clknet_leaf_213_clk),
    .Q(\register_file[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15893_ (.D(_00281_),
    .CLK(clknet_leaf_216_clk),
    .Q(\register_file[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15894_ (.D(_00282_),
    .CLK(clknet_leaf_203_clk),
    .Q(\register_file[11][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15895_ (.D(_00283_),
    .CLK(clknet_leaf_217_clk),
    .Q(\register_file[11][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15896_ (.D(_00284_),
    .CLK(clknet_leaf_264_clk),
    .Q(\register_file[11][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15897_ (.D(_00285_),
    .CLK(clknet_leaf_261_clk),
    .Q(\register_file[11][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15898_ (.D(_00286_),
    .CLK(clknet_leaf_265_clk),
    .Q(\register_file[11][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15899_ (.D(_00287_),
    .CLK(clknet_leaf_265_clk),
    .Q(\register_file[11][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15900_ (.D(_00288_),
    .CLK(clknet_leaf_283_clk),
    .Q(\register_file[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15901_ (.D(_00289_),
    .CLK(clknet_leaf_280_clk),
    .Q(\register_file[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15902_ (.D(_00290_),
    .CLK(clknet_leaf_303_clk),
    .Q(\register_file[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15903_ (.D(_00291_),
    .CLK(clknet_leaf_10_clk),
    .Q(\register_file[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15904_ (.D(_00292_),
    .CLK(clknet_leaf_7_clk),
    .Q(\register_file[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15905_ (.D(_00293_),
    .CLK(clknet_leaf_23_clk),
    .Q(\register_file[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15906_ (.D(_00294_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(\register_file[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15907_ (.D(_00295_),
    .CLK(clknet_leaf_50_clk),
    .Q(\register_file[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15908_ (.D(_00296_),
    .CLK(clknet_leaf_62_clk),
    .Q(\register_file[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15909_ (.D(_00297_),
    .CLK(clknet_leaf_63_clk),
    .Q(\register_file[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15910_ (.D(_00298_),
    .CLK(clknet_leaf_109_clk),
    .Q(\register_file[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15911_ (.D(_00299_),
    .CLK(clknet_leaf_109_clk),
    .Q(\register_file[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15912_ (.D(_00300_),
    .CLK(clknet_leaf_109_clk),
    .Q(\register_file[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15913_ (.D(_00301_),
    .CLK(clknet_leaf_111_clk),
    .Q(\register_file[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15914_ (.D(_00302_),
    .CLK(clknet_leaf_112_clk),
    .Q(\register_file[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15915_ (.D(_00303_),
    .CLK(clknet_leaf_112_clk),
    .Q(\register_file[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15916_ (.D(_00304_),
    .CLK(clknet_leaf_122_clk),
    .Q(\register_file[10][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15917_ (.D(_00305_),
    .CLK(clknet_leaf_121_clk),
    .Q(\register_file[10][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15918_ (.D(_00306_),
    .CLK(clknet_leaf_187_clk),
    .Q(\register_file[10][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15919_ (.D(_00307_),
    .CLK(clknet_leaf_186_clk),
    .Q(\register_file[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15920_ (.D(_00308_),
    .CLK(clknet_leaf_186_clk),
    .Q(\register_file[10][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15921_ (.D(_00309_),
    .CLK(clknet_leaf_185_clk),
    .Q(\register_file[10][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15922_ (.D(_00310_),
    .CLK(clknet_leaf_185_clk),
    .Q(\register_file[10][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15923_ (.D(_00311_),
    .CLK(clknet_leaf_213_clk),
    .Q(\register_file[10][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15924_ (.D(_00312_),
    .CLK(clknet_leaf_209_clk),
    .Q(\register_file[10][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15925_ (.D(_00313_),
    .CLK(clknet_leaf_218_clk),
    .Q(\register_file[10][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15926_ (.D(_00314_),
    .CLK(clknet_leaf_203_clk),
    .Q(\register_file[10][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15927_ (.D(_00315_),
    .CLK(clknet_leaf_220_clk),
    .Q(\register_file[10][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15928_ (.D(_00316_),
    .CLK(clknet_leaf_264_clk),
    .Q(\register_file[10][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15929_ (.D(_00317_),
    .CLK(clknet_leaf_256_clk),
    .Q(\register_file[10][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15930_ (.D(_00318_),
    .CLK(clknet_leaf_256_clk),
    .Q(\register_file[10][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15931_ (.D(_00319_),
    .CLK(clknet_leaf_265_clk),
    .Q(\register_file[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15932_ (.D(_00320_),
    .CLK(clknet_leaf_287_clk),
    .Q(\register_file[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15933_ (.D(_00321_),
    .CLK(clknet_leaf_307_clk),
    .Q(\register_file[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15934_ (.D(_00322_),
    .CLK(clknet_leaf_305_clk),
    .Q(\register_file[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15935_ (.D(_00323_),
    .CLK(clknet_leaf_3_clk),
    .Q(\register_file[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15936_ (.D(_00324_),
    .CLK(clknet_leaf_2_clk),
    .Q(\register_file[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15937_ (.D(_00325_),
    .CLK(clknet_leaf_4_clk),
    .Q(\register_file[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15938_ (.D(_00326_),
    .CLK(clknet_leaf_4_clk),
    .Q(\register_file[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15939_ (.D(_00327_),
    .CLK(clknet_leaf_14_clk),
    .Q(\register_file[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15940_ (.D(_00328_),
    .CLK(clknet_leaf_58_clk),
    .Q(\register_file[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15941_ (.D(_00329_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\register_file[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15942_ (.D(_00330_),
    .CLK(clknet_leaf_49_clk),
    .Q(\register_file[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15943_ (.D(_00331_),
    .CLK(clknet_leaf_43_clk),
    .Q(\register_file[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15944_ (.D(_00332_),
    .CLK(clknet_leaf_44_clk),
    .Q(\register_file[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15945_ (.D(_00333_),
    .CLK(clknet_leaf_41_clk),
    .Q(\register_file[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15946_ (.D(_00334_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\register_file[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15947_ (.D(_00335_),
    .CLK(clknet_leaf_115_clk),
    .Q(\register_file[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15948_ (.D(_00336_),
    .CLK(clknet_leaf_117_clk),
    .Q(\register_file[8][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15949_ (.D(_00337_),
    .CLK(clknet_leaf_117_clk),
    .Q(\register_file[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15950_ (.D(_00338_),
    .CLK(clknet_leaf_189_clk),
    .Q(\register_file[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15951_ (.D(_00339_),
    .CLK(clknet_leaf_189_clk),
    .Q(\register_file[8][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15952_ (.D(_00340_),
    .CLK(clknet_leaf_216_clk),
    .Q(\register_file[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15953_ (.D(_00341_),
    .CLK(clknet_leaf_216_clk),
    .Q(\register_file[8][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15954_ (.D(_00342_),
    .CLK(clknet_leaf_216_clk),
    .Q(\register_file[8][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15955_ (.D(_00343_),
    .CLK(clknet_leaf_226_clk),
    .Q(\register_file[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15956_ (.D(_00344_),
    .CLK(clknet_leaf_221_clk),
    .Q(\register_file[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15957_ (.D(_00345_),
    .CLK(clknet_leaf_221_clk),
    .Q(\register_file[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15958_ (.D(_00346_),
    .CLK(clknet_leaf_239_clk),
    .Q(\register_file[8][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15959_ (.D(_00347_),
    .CLK(clknet_leaf_239_clk),
    .Q(\register_file[8][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15960_ (.D(_00348_),
    .CLK(clknet_leaf_242_clk),
    .Q(\register_file[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15961_ (.D(_00349_),
    .CLK(clknet_leaf_257_clk),
    .Q(\register_file[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15962_ (.D(_00350_),
    .CLK(clknet_leaf_253_clk),
    .Q(\register_file[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15963_ (.D(_00351_),
    .CLK(clknet_leaf_285_clk),
    .Q(\register_file[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15964_ (.D(_00352_),
    .CLK(clknet_leaf_293_clk),
    .Q(\register_file[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15965_ (.D(_00353_),
    .CLK(clknet_leaf_307_clk),
    .Q(\register_file[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15966_ (.D(_00354_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\register_file[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15967_ (.D(_00355_),
    .CLK(clknet_leaf_1_clk),
    .Q(\register_file[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15968_ (.D(_00356_),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\register_file[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15969_ (.D(_00357_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15970_ (.D(_00358_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15971_ (.D(_00359_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15972_ (.D(_00360_),
    .CLK(clknet_leaf_313_clk),
    .Q(\register_file[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15973_ (.D(_00361_),
    .CLK(clknet_leaf_313_clk),
    .Q(\register_file[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15974_ (.D(_00362_),
    .CLK(clknet_leaf_309_clk),
    .Q(\register_file[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15975_ (.D(_00363_),
    .CLK(clknet_leaf_297_clk),
    .Q(\register_file[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15976_ (.D(_00364_),
    .CLK(clknet_leaf_297_clk),
    .Q(\register_file[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15977_ (.D(_00365_),
    .CLK(clknet_leaf_291_clk),
    .Q(\register_file[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15978_ (.D(_00366_),
    .CLK(clknet_leaf_291_clk),
    .Q(\register_file[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15979_ (.D(_00367_),
    .CLK(clknet_leaf_250_clk),
    .Q(\register_file[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15980_ (.D(_00368_),
    .CLK(clknet_leaf_249_clk),
    .Q(\register_file[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15981_ (.D(_00369_),
    .CLK(clknet_leaf_247_clk),
    .Q(\register_file[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15982_ (.D(_00370_),
    .CLK(clknet_leaf_245_clk),
    .Q(\register_file[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15983_ (.D(_00371_),
    .CLK(clknet_leaf_245_clk),
    .Q(\register_file[7][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15984_ (.D(_00372_),
    .CLK(clknet_leaf_230_clk),
    .Q(\register_file[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15985_ (.D(_00373_),
    .CLK(clknet_leaf_229_clk),
    .Q(\register_file[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15986_ (.D(_00374_),
    .CLK(clknet_leaf_229_clk),
    .Q(\register_file[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15987_ (.D(_00375_),
    .CLK(clknet_leaf_228_clk),
    .Q(\register_file[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15988_ (.D(_00376_),
    .CLK(clknet_leaf_229_clk),
    .Q(\register_file[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15989_ (.D(_00377_),
    .CLK(clknet_leaf_233_clk),
    .Q(\register_file[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15990_ (.D(_00378_),
    .CLK(clknet_leaf_237_clk),
    .Q(\register_file[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15991_ (.D(_00379_),
    .CLK(clknet_leaf_235_clk),
    .Q(\register_file[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15992_ (.D(_00380_),
    .CLK(clknet_leaf_244_clk),
    .Q(\register_file[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15993_ (.D(_00381_),
    .CLK(clknet_leaf_243_clk),
    .Q(\register_file[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15994_ (.D(_00382_),
    .CLK(clknet_leaf_252_clk),
    .Q(\register_file[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15995_ (.D(_00383_),
    .CLK(clknet_leaf_288_clk),
    .Q(\register_file[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15996_ (.D(_00384_),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\register_file[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15997_ (.D(_00385_),
    .CLK(clknet_leaf_307_clk),
    .Q(\register_file[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15998_ (.D(_00386_),
    .CLK(clknet_leaf_306_clk),
    .Q(\register_file[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15999_ (.D(_00387_),
    .CLK(clknet_leaf_0_clk),
    .Q(\register_file[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16000_ (.D(_00388_),
    .CLK(clknet_leaf_0_clk),
    .Q(\register_file[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16001_ (.D(_00389_),
    .CLK(clknet_leaf_0_clk),
    .Q(\register_file[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16002_ (.D(_00390_),
    .CLK(clknet_leaf_0_clk),
    .Q(\register_file[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16003_ (.D(_00391_),
    .CLK(clknet_leaf_0_clk),
    .Q(\register_file[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16004_ (.D(_00392_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16005_ (.D(_00393_),
    .CLK(clknet_leaf_313_clk),
    .Q(\register_file[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16006_ (.D(_00394_),
    .CLK(clknet_leaf_309_clk),
    .Q(\register_file[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16007_ (.D(_00395_),
    .CLK(clknet_leaf_297_clk),
    .Q(\register_file[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16008_ (.D(_00396_),
    .CLK(clknet_leaf_296_clk),
    .Q(\register_file[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16009_ (.D(_00397_),
    .CLK(clknet_leaf_292_clk),
    .Q(\register_file[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16010_ (.D(_00398_),
    .CLK(clknet_leaf_292_clk),
    .Q(\register_file[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16011_ (.D(_00399_),
    .CLK(clknet_leaf_250_clk),
    .Q(\register_file[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16012_ (.D(_00400_),
    .CLK(clknet_leaf_249_clk),
    .Q(\register_file[6][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16013_ (.D(_00401_),
    .CLK(clknet_leaf_247_clk),
    .Q(\register_file[6][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16014_ (.D(_00402_),
    .CLK(clknet_leaf_246_clk),
    .Q(\register_file[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16015_ (.D(_00403_),
    .CLK(clknet_leaf_244_clk),
    .Q(\register_file[6][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16016_ (.D(_00404_),
    .CLK(clknet_leaf_229_clk),
    .Q(\register_file[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16017_ (.D(_00405_),
    .CLK(clknet_leaf_229_clk),
    .Q(\register_file[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16018_ (.D(_00406_),
    .CLK(clknet_leaf_229_clk),
    .Q(\register_file[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16019_ (.D(_00407_),
    .CLK(clknet_leaf_228_clk),
    .Q(\register_file[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16020_ (.D(_00408_),
    .CLK(clknet_leaf_228_clk),
    .Q(\register_file[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16021_ (.D(_00409_),
    .CLK(clknet_leaf_238_clk),
    .Q(\register_file[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16022_ (.D(_00410_),
    .CLK(clknet_leaf_237_clk),
    .Q(\register_file[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16023_ (.D(_00411_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\register_file[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16024_ (.D(_00412_),
    .CLK(clknet_leaf_243_clk),
    .Q(\register_file[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16025_ (.D(_00413_),
    .CLK(clknet_leaf_243_clk),
    .Q(\register_file[6][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16026_ (.D(_00414_),
    .CLK(clknet_leaf_252_clk),
    .Q(\register_file[6][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16027_ (.D(_00415_),
    .CLK(clknet_leaf_252_clk),
    .Q(\register_file[6][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16028_ (.D(_00416_),
    .CLK(clknet_leaf_293_clk),
    .Q(\register_file[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16029_ (.D(_00417_),
    .CLK(clknet_leaf_298_clk),
    .Q(\register_file[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16030_ (.D(_00418_),
    .CLK(clknet_leaf_298_clk),
    .Q(\register_file[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16031_ (.D(_00419_),
    .CLK(clknet_leaf_0_clk),
    .Q(\register_file[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16032_ (.D(_00420_),
    .CLK(clknet_leaf_1_clk),
    .Q(\register_file[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16033_ (.D(_00421_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16034_ (.D(_00422_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16035_ (.D(_00423_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16036_ (.D(_00424_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16037_ (.D(_00425_),
    .CLK(clknet_leaf_314_clk),
    .Q(\register_file[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16038_ (.D(_00426_),
    .CLK(clknet_leaf_309_clk),
    .Q(\register_file[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16039_ (.D(_00427_),
    .CLK(clknet_leaf_296_clk),
    .Q(\register_file[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16040_ (.D(_00428_),
    .CLK(clknet_leaf_296_clk),
    .Q(\register_file[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16041_ (.D(_00429_),
    .CLK(clknet_leaf_291_clk),
    .Q(\register_file[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16042_ (.D(_00430_),
    .CLK(clknet_leaf_289_clk),
    .Q(\register_file[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16043_ (.D(_00431_),
    .CLK(clknet_leaf_289_clk),
    .Q(\register_file[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16044_ (.D(_00432_),
    .CLK(clknet_leaf_251_clk),
    .Q(\register_file[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16045_ (.D(_00433_),
    .CLK(clknet_leaf_249_clk),
    .Q(\register_file[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16046_ (.D(_00434_),
    .CLK(clknet_leaf_245_clk),
    .Q(\register_file[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16047_ (.D(_00435_),
    .CLK(clknet_leaf_245_clk),
    .Q(\register_file[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16048_ (.D(_00436_),
    .CLK(clknet_leaf_230_clk),
    .Q(\register_file[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16049_ (.D(_00437_),
    .CLK(clknet_leaf_230_clk),
    .Q(\register_file[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16050_ (.D(_00438_),
    .CLK(clknet_leaf_230_clk),
    .Q(\register_file[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16051_ (.D(_00439_),
    .CLK(clknet_leaf_231_clk),
    .Q(\register_file[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16052_ (.D(_00440_),
    .CLK(clknet_leaf_230_clk),
    .Q(\register_file[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16053_ (.D(_00441_),
    .CLK(clknet_leaf_233_clk),
    .Q(\register_file[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16054_ (.D(_00442_),
    .CLK(clknet_leaf_234_clk),
    .Q(\register_file[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16055_ (.D(_00443_),
    .CLK(clknet_leaf_235_clk),
    .Q(\register_file[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16056_ (.D(_00444_),
    .CLK(clknet_leaf_244_clk),
    .Q(\register_file[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16057_ (.D(_00445_),
    .CLK(clknet_leaf_242_clk),
    .Q(\register_file[5][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16058_ (.D(_00446_),
    .CLK(clknet_leaf_248_clk),
    .Q(\register_file[5][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16059_ (.D(_00447_),
    .CLK(clknet_leaf_288_clk),
    .Q(\register_file[5][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16060_ (.D(_00448_),
    .CLK(clknet_leaf_293_clk),
    .Q(\register_file[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16061_ (.D(_00449_),
    .CLK(clknet_leaf_300_clk),
    .Q(\register_file[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16062_ (.D(_00450_),
    .CLK(clknet_leaf_300_clk),
    .Q(\register_file[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16063_ (.D(_00451_),
    .CLK(clknet_leaf_306_clk),
    .Q(\register_file[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16064_ (.D(_00452_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\register_file[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16065_ (.D(_00453_),
    .CLK(clknet_leaf_313_clk),
    .Q(\register_file[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16066_ (.D(_00454_),
    .CLK(clknet_leaf_310_clk),
    .Q(\register_file[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16067_ (.D(_00455_),
    .CLK(clknet_leaf_310_clk),
    .Q(\register_file[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16068_ (.D(_00456_),
    .CLK(clknet_leaf_313_clk),
    .Q(\register_file[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16069_ (.D(_00457_),
    .CLK(clknet_leaf_310_clk),
    .Q(\register_file[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16070_ (.D(_00458_),
    .CLK(clknet_leaf_309_clk),
    .Q(\register_file[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16071_ (.D(_00459_),
    .CLK(clknet_leaf_295_clk),
    .Q(\register_file[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16072_ (.D(_00460_),
    .CLK(clknet_leaf_295_clk),
    .Q(\register_file[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16073_ (.D(_00461_),
    .CLK(clknet_leaf_289_clk),
    .Q(\register_file[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16074_ (.D(_00462_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\register_file[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16075_ (.D(_00463_),
    .CLK(clknet_leaf_251_clk),
    .Q(\register_file[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16076_ (.D(_00464_),
    .CLK(clknet_leaf_251_clk),
    .Q(\register_file[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16077_ (.D(_00465_),
    .CLK(clknet_leaf_247_clk),
    .Q(\register_file[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16078_ (.D(_00466_),
    .CLK(clknet_leaf_246_clk),
    .Q(\register_file[4][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16079_ (.D(_00467_),
    .CLK(clknet_leaf_234_clk),
    .Q(\register_file[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16080_ (.D(_00468_),
    .CLK(clknet_leaf_234_clk),
    .Q(\register_file[4][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16081_ (.D(_00469_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(\register_file[4][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16082_ (.D(_00470_),
    .CLK(clknet_leaf_231_clk),
    .Q(\register_file[4][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16083_ (.D(_00471_),
    .CLK(clknet_leaf_231_clk),
    .Q(\register_file[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16084_ (.D(_00472_),
    .CLK(clknet_leaf_230_clk),
    .Q(\register_file[4][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16085_ (.D(_00473_),
    .CLK(clknet_leaf_233_clk),
    .Q(\register_file[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16086_ (.D(_00474_),
    .CLK(clknet_leaf_234_clk),
    .Q(\register_file[4][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16087_ (.D(_00475_),
    .CLK(clknet_leaf_234_clk),
    .Q(\register_file[4][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16088_ (.D(_00476_),
    .CLK(clknet_leaf_235_clk),
    .Q(\register_file[4][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16089_ (.D(_00477_),
    .CLK(clknet_leaf_248_clk),
    .Q(\register_file[4][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16090_ (.D(_00478_),
    .CLK(clknet_leaf_248_clk),
    .Q(\register_file[4][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16091_ (.D(_00479_),
    .CLK(clknet_leaf_288_clk),
    .Q(\register_file[4][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16092_ (.D(_00480_),
    .CLK(clknet_leaf_301_clk),
    .Q(\register_file[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16093_ (.D(_00481_),
    .CLK(clknet_leaf_299_clk),
    .Q(\register_file[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16094_ (.D(_00482_),
    .CLK(clknet_leaf_299_clk),
    .Q(\register_file[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16095_ (.D(_00483_),
    .CLK(clknet_leaf_3_clk),
    .Q(\register_file[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16096_ (.D(_00484_),
    .CLK(clknet_leaf_3_clk),
    .Q(\register_file[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16097_ (.D(_00485_),
    .CLK(clknet_leaf_14_clk),
    .Q(\register_file[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16098_ (.D(_00486_),
    .CLK(clknet_leaf_14_clk),
    .Q(\register_file[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16099_ (.D(_00487_),
    .CLK(clknet_leaf_14_clk),
    .Q(\register_file[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16100_ (.D(_00488_),
    .CLK(clknet_leaf_54_clk),
    .Q(\register_file[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16101_ (.D(_00489_),
    .CLK(clknet_leaf_54_clk),
    .Q(\register_file[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16102_ (.D(_00490_),
    .CLK(clknet_leaf_44_clk),
    .Q(\register_file[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16103_ (.D(_00491_),
    .CLK(clknet_leaf_42_clk),
    .Q(\register_file[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16104_ (.D(_00492_),
    .CLK(clknet_leaf_42_clk),
    .Q(\register_file[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16105_ (.D(_00493_),
    .CLK(clknet_leaf_41_clk),
    .Q(\register_file[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16106_ (.D(_00494_),
    .CLK(clknet_leaf_41_clk),
    .Q(\register_file[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16107_ (.D(_00495_),
    .CLK(clknet_leaf_193_clk),
    .Q(\register_file[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16108_ (.D(_00496_),
    .CLK(clknet_leaf_193_clk),
    .Q(\register_file[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16109_ (.D(_00497_),
    .CLK(clknet_leaf_192_clk),
    .Q(\register_file[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16110_ (.D(_00498_),
    .CLK(clknet_leaf_192_clk),
    .Q(\register_file[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16111_ (.D(_00499_),
    .CLK(clknet_leaf_190_clk),
    .Q(\register_file[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16112_ (.D(_00500_),
    .CLK(clknet_leaf_226_clk),
    .Q(\register_file[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16113_ (.D(_00501_),
    .CLK(clknet_leaf_226_clk),
    .Q(\register_file[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16114_ (.D(_00502_),
    .CLK(clknet_leaf_229_clk),
    .Q(\register_file[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16115_ (.D(_00503_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(\register_file[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16116_ (.D(_00504_),
    .CLK(clknet_leaf_221_clk),
    .Q(\register_file[3][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16117_ (.D(_00505_),
    .CLK(clknet_leaf_221_clk),
    .Q(\register_file[3][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16118_ (.D(_00506_),
    .CLK(clknet_leaf_238_clk),
    .Q(\register_file[3][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16119_ (.D(_00507_),
    .CLK(clknet_leaf_239_clk),
    .Q(\register_file[3][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16120_ (.D(_00508_),
    .CLK(clknet_leaf_241_clk),
    .Q(\register_file[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16121_ (.D(_00509_),
    .CLK(clknet_leaf_241_clk),
    .Q(\register_file[3][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16122_ (.D(_00510_),
    .CLK(clknet_leaf_253_clk),
    .Q(\register_file[3][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16123_ (.D(_00511_),
    .CLK(clknet_leaf_288_clk),
    .Q(\register_file[3][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16124_ (.D(_00512_),
    .CLK(clknet_leaf_37_clk),
    .Q(\register_file[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16125_ (.D(_00513_),
    .CLK(clknet_leaf_34_clk),
    .Q(\register_file[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16126_ (.D(_00514_),
    .CLK(clknet_leaf_33_clk),
    .Q(\register_file[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16127_ (.D(_00515_),
    .CLK(clknet_leaf_18_clk),
    .Q(\register_file[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16128_ (.D(_00516_),
    .CLK(clknet_leaf_18_clk),
    .Q(\register_file[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16129_ (.D(_00517_),
    .CLK(clknet_leaf_67_clk),
    .Q(\register_file[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16130_ (.D(_00518_),
    .CLK(clknet_leaf_60_clk),
    .Q(\register_file[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16131_ (.D(_00519_),
    .CLK(clknet_leaf_61_clk),
    .Q(\register_file[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16132_ (.D(_00520_),
    .CLK(clknet_leaf_76_clk),
    .Q(\register_file[31][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16133_ (.D(_00521_),
    .CLK(clknet_leaf_79_clk),
    .Q(\register_file[31][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16134_ (.D(_00522_),
    .CLK(clknet_leaf_90_clk),
    .Q(\register_file[31][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16135_ (.D(_00523_),
    .CLK(clknet_leaf_92_clk),
    .Q(\register_file[31][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16136_ (.D(_00524_),
    .CLK(clknet_leaf_90_clk),
    .Q(\register_file[31][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16137_ (.D(_00525_),
    .CLK(clknet_leaf_95_clk),
    .Q(\register_file[31][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16138_ (.D(_00526_),
    .CLK(clknet_leaf_93_clk),
    .Q(\register_file[31][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16139_ (.D(_00527_),
    .CLK(clknet_leaf_98_clk),
    .Q(\register_file[31][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16140_ (.D(_00528_),
    .CLK(clknet_leaf_139_clk),
    .Q(\register_file[31][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16141_ (.D(_00529_),
    .CLK(clknet_leaf_140_clk),
    .Q(\register_file[31][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16142_ (.D(_00530_),
    .CLK(clknet_leaf_153_clk),
    .Q(\register_file[31][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16143_ (.D(_00531_),
    .CLK(clknet_leaf_153_clk),
    .Q(\register_file[31][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16144_ (.D(_00532_),
    .CLK(clknet_leaf_156_clk),
    .Q(\register_file[31][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16145_ (.D(_00533_),
    .CLK(clknet_leaf_156_clk),
    .Q(\register_file[31][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16146_ (.D(_00534_),
    .CLK(clknet_leaf_156_clk),
    .Q(\register_file[31][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16147_ (.D(_00535_),
    .CLK(clknet_leaf_151_clk),
    .Q(\register_file[31][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16148_ (.D(_00536_),
    .CLK(clknet_leaf_151_clk),
    .Q(\register_file[31][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16149_ (.D(_00537_),
    .CLK(clknet_leaf_181_clk),
    .Q(\register_file[31][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16150_ (.D(_00538_),
    .CLK(clknet_leaf_181_clk),
    .Q(\register_file[31][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16151_ (.D(_00539_),
    .CLK(clknet_leaf_190_clk),
    .Q(\register_file[31][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16152_ (.D(_00540_),
    .CLK(clknet_leaf_190_clk),
    .Q(\register_file[31][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16153_ (.D(_00541_),
    .CLK(clknet_leaf_191_clk),
    .Q(\register_file[31][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16154_ (.D(_00542_),
    .CLK(clknet_leaf_269_clk),
    .Q(\register_file[31][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16155_ (.D(_00543_),
    .CLK(clknet_leaf_39_clk),
    .Q(\register_file[31][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16156_ (.D(_00544_),
    .CLK(clknet_leaf_35_clk),
    .Q(\register_file[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16157_ (.D(_00545_),
    .CLK(clknet_leaf_35_clk),
    .Q(\register_file[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16158_ (.D(_00546_),
    .CLK(clknet_leaf_24_clk),
    .Q(\register_file[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16159_ (.D(_00547_),
    .CLK(clknet_leaf_17_clk),
    .Q(\register_file[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16160_ (.D(_00548_),
    .CLK(clknet_leaf_12_clk),
    .Q(\register_file[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16161_ (.D(_00549_),
    .CLK(clknet_leaf_65_clk),
    .Q(\register_file[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16162_ (.D(_00550_),
    .CLK(clknet_leaf_65_clk),
    .Q(\register_file[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16163_ (.D(_00551_),
    .CLK(clknet_leaf_65_clk),
    .Q(\register_file[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16164_ (.D(_00552_),
    .CLK(clknet_leaf_75_clk),
    .Q(\register_file[25][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16165_ (.D(_00553_),
    .CLK(clknet_leaf_80_clk),
    .Q(\register_file[25][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16166_ (.D(_00554_),
    .CLK(clknet_leaf_91_clk),
    .Q(\register_file[25][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16167_ (.D(_00555_),
    .CLK(clknet_leaf_92_clk),
    .Q(\register_file[25][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16168_ (.D(_00556_),
    .CLK(clknet_leaf_92_clk),
    .Q(\register_file[25][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16169_ (.D(_00557_),
    .CLK(clknet_leaf_93_clk),
    .Q(\register_file[25][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16170_ (.D(_00558_),
    .CLK(clknet_leaf_93_clk),
    .Q(\register_file[25][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16171_ (.D(_00559_),
    .CLK(clknet_leaf_98_clk),
    .Q(\register_file[25][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16172_ (.D(_00560_),
    .CLK(clknet_leaf_138_clk),
    .Q(\register_file[25][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16173_ (.D(_00561_),
    .CLK(clknet_leaf_138_clk),
    .Q(\register_file[25][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16174_ (.D(_00562_),
    .CLK(clknet_leaf_143_clk),
    .Q(\register_file[25][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16175_ (.D(_00563_),
    .CLK(clknet_leaf_144_clk),
    .Q(\register_file[25][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16176_ (.D(_00564_),
    .CLK(clknet_leaf_154_clk),
    .Q(\register_file[25][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16177_ (.D(_00565_),
    .CLK(clknet_leaf_155_clk),
    .Q(\register_file[25][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16178_ (.D(_00566_),
    .CLK(clknet_leaf_155_clk),
    .Q(\register_file[25][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16179_ (.D(_00567_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\register_file[25][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16180_ (.D(_00568_),
    .CLK(clknet_leaf_162_clk),
    .Q(\register_file[25][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16181_ (.D(_00569_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(\register_file[25][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16182_ (.D(_00570_),
    .CLK(clknet_leaf_182_clk),
    .Q(\register_file[25][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16183_ (.D(_00571_),
    .CLK(clknet_leaf_190_clk),
    .Q(\register_file[25][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16184_ (.D(_00572_),
    .CLK(clknet_leaf_191_clk),
    .Q(\register_file[25][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16185_ (.D(_00573_),
    .CLK(clknet_leaf_196_clk),
    .Q(\register_file[25][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16186_ (.D(_00574_),
    .CLK(clknet_leaf_40_clk),
    .Q(\register_file[25][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16187_ (.D(_00575_),
    .CLK(clknet_leaf_40_clk),
    .Q(\register_file[25][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16188_ (.D(_00576_),
    .CLK(clknet_leaf_35_clk),
    .Q(\register_file[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16189_ (.D(_00577_),
    .CLK(clknet_leaf_34_clk),
    .Q(\register_file[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16190_ (.D(_00578_),
    .CLK(clknet_leaf_33_clk),
    .Q(\register_file[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16191_ (.D(_00579_),
    .CLK(clknet_leaf_11_clk),
    .Q(\register_file[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16192_ (.D(_00580_),
    .CLK(clknet_leaf_11_clk),
    .Q(\register_file[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16193_ (.D(_00581_),
    .CLK(clknet_leaf_70_clk),
    .Q(\register_file[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16194_ (.D(_00582_),
    .CLK(clknet_leaf_70_clk),
    .Q(\register_file[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16195_ (.D(_00583_),
    .CLK(clknet_leaf_71_clk),
    .Q(\register_file[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16196_ (.D(_00584_),
    .CLK(clknet_leaf_76_clk),
    .Q(\register_file[24][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16197_ (.D(_00585_),
    .CLK(clknet_leaf_80_clk),
    .Q(\register_file[24][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16198_ (.D(_00586_),
    .CLK(clknet_leaf_91_clk),
    .Q(\register_file[24][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16199_ (.D(_00587_),
    .CLK(clknet_leaf_92_clk),
    .Q(\register_file[24][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16200_ (.D(_00588_),
    .CLK(clknet_leaf_92_clk),
    .Q(\register_file[24][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16201_ (.D(_00589_),
    .CLK(clknet_leaf_96_clk),
    .Q(\register_file[24][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16202_ (.D(_00590_),
    .CLK(clknet_leaf_96_clk),
    .Q(\register_file[24][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16203_ (.D(_00591_),
    .CLK(clknet_leaf_97_clk),
    .Q(\register_file[24][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16204_ (.D(_00592_),
    .CLK(clknet_leaf_98_clk),
    .Q(\register_file[24][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16205_ (.D(_00593_),
    .CLK(clknet_leaf_138_clk),
    .Q(\register_file[24][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16206_ (.D(_00594_),
    .CLK(clknet_leaf_143_clk),
    .Q(\register_file[24][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16207_ (.D(_00595_),
    .CLK(clknet_leaf_143_clk),
    .Q(\register_file[24][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16208_ (.D(_00596_),
    .CLK(clknet_leaf_154_clk),
    .Q(\register_file[24][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16209_ (.D(_00597_),
    .CLK(clknet_leaf_155_clk),
    .Q(\register_file[24][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16210_ (.D(_00598_),
    .CLK(clknet_leaf_155_clk),
    .Q(\register_file[24][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16211_ (.D(_00599_),
    .CLK(clknet_leaf_157_clk),
    .Q(\register_file[24][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16212_ (.D(_00600_),
    .CLK(clknet_leaf_157_clk),
    .Q(\register_file[24][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16213_ (.D(_00601_),
    .CLK(clknet_leaf_183_clk),
    .Q(\register_file[24][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16214_ (.D(_00602_),
    .CLK(clknet_leaf_207_clk),
    .Q(\register_file[24][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16215_ (.D(_00603_),
    .CLK(clknet_leaf_197_clk),
    .Q(\register_file[24][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16216_ (.D(_00604_),
    .CLK(clknet_leaf_196_clk),
    .Q(\register_file[24][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16217_ (.D(_00605_),
    .CLK(clknet_leaf_196_clk),
    .Q(\register_file[24][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16218_ (.D(_00606_),
    .CLK(clknet_leaf_38_clk),
    .Q(\register_file[24][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16219_ (.D(_00607_),
    .CLK(clknet_leaf_39_clk),
    .Q(\register_file[24][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16220_ (.D(_00608_),
    .CLK(clknet_leaf_38_clk),
    .Q(\register_file[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16221_ (.D(_00609_),
    .CLK(clknet_leaf_34_clk),
    .Q(\register_file[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16222_ (.D(_00610_),
    .CLK(clknet_leaf_33_clk),
    .Q(\register_file[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16223_ (.D(_00611_),
    .CLK(clknet_leaf_24_clk),
    .Q(\register_file[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16224_ (.D(_00612_),
    .CLK(clknet_leaf_23_clk),
    .Q(\register_file[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16225_ (.D(_00613_),
    .CLK(clknet_leaf_72_clk),
    .Q(\register_file[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16226_ (.D(_00614_),
    .CLK(clknet_leaf_72_clk),
    .Q(\register_file[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16227_ (.D(_00615_),
    .CLK(clknet_leaf_78_clk),
    .Q(\register_file[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16228_ (.D(_00616_),
    .CLK(clknet_leaf_77_clk),
    .Q(\register_file[23][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16229_ (.D(_00617_),
    .CLK(clknet_leaf_78_clk),
    .Q(\register_file[23][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16230_ (.D(_00618_),
    .CLK(clknet_leaf_82_clk),
    .Q(\register_file[23][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16231_ (.D(_00619_),
    .CLK(clknet_leaf_90_clk),
    .Q(\register_file[23][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16232_ (.D(_00620_),
    .CLK(clknet_leaf_93_clk),
    .Q(\register_file[23][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16233_ (.D(_00621_),
    .CLK(clknet_leaf_95_clk),
    .Q(\register_file[23][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16234_ (.D(_00622_),
    .CLK(clknet_leaf_97_clk),
    .Q(\register_file[23][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16235_ (.D(_00623_),
    .CLK(clknet_leaf_136_clk),
    .Q(\register_file[23][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16236_ (.D(_00624_),
    .CLK(clknet_leaf_137_clk),
    .Q(\register_file[23][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16237_ (.D(_00625_),
    .CLK(clknet_leaf_139_clk),
    .Q(\register_file[23][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16238_ (.D(_00626_),
    .CLK(clknet_leaf_145_clk),
    .Q(\register_file[23][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16239_ (.D(_00627_),
    .CLK(clknet_leaf_153_clk),
    .Q(\register_file[23][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16240_ (.D(_00628_),
    .CLK(clknet_leaf_151_clk),
    .Q(\register_file[23][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16241_ (.D(_00629_),
    .CLK(clknet_leaf_156_clk),
    .Q(\register_file[23][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16242_ (.D(_00630_),
    .CLK(clknet_leaf_156_clk),
    .Q(\register_file[23][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16243_ (.D(_00631_),
    .CLK(clknet_leaf_181_clk),
    .Q(\register_file[23][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16244_ (.D(_00632_),
    .CLK(clknet_leaf_181_clk),
    .Q(\register_file[23][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16245_ (.D(_00633_),
    .CLK(clknet_leaf_183_clk),
    .Q(\register_file[23][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16246_ (.D(_00634_),
    .CLK(clknet_leaf_183_clk),
    .Q(\register_file[23][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16247_ (.D(_00635_),
    .CLK(clknet_leaf_190_clk),
    .Q(\register_file[23][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16248_ (.D(_00636_),
    .CLK(clknet_leaf_193_clk),
    .Q(\register_file[23][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16249_ (.D(_00637_),
    .CLK(clknet_leaf_193_clk),
    .Q(\register_file[23][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16250_ (.D(_00638_),
    .CLK(clknet_leaf_269_clk),
    .Q(\register_file[23][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16251_ (.D(_00639_),
    .CLK(clknet_leaf_269_clk),
    .Q(\register_file[23][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16252_ (.D(_00640_),
    .CLK(clknet_leaf_38_clk),
    .Q(\register_file[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16253_ (.D(_00641_),
    .CLK(clknet_leaf_34_clk),
    .Q(\register_file[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16254_ (.D(_00642_),
    .CLK(clknet_leaf_43_clk),
    .Q(\register_file[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16255_ (.D(_00643_),
    .CLK(clknet_leaf_24_clk),
    .Q(\register_file[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16256_ (.D(_00644_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\register_file[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16257_ (.D(_00645_),
    .CLK(clknet_leaf_71_clk),
    .Q(\register_file[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16258_ (.D(_00646_),
    .CLK(clknet_leaf_71_clk),
    .Q(\register_file[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16259_ (.D(_00647_),
    .CLK(clknet_leaf_78_clk),
    .Q(\register_file[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16260_ (.D(_00648_),
    .CLK(clknet_leaf_75_clk),
    .Q(\register_file[22][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16261_ (.D(_00649_),
    .CLK(clknet_leaf_75_clk),
    .Q(\register_file[22][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16262_ (.D(_00650_),
    .CLK(clknet_leaf_91_clk),
    .Q(\register_file[22][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16263_ (.D(_00651_),
    .CLK(clknet_leaf_91_clk),
    .Q(\register_file[22][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16264_ (.D(_00652_),
    .CLK(clknet_leaf_91_clk),
    .Q(\register_file[22][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16265_ (.D(_00653_),
    .CLK(clknet_leaf_96_clk),
    .Q(\register_file[22][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16266_ (.D(_00654_),
    .CLK(clknet_leaf_96_clk),
    .Q(\register_file[22][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16267_ (.D(_00655_),
    .CLK(clknet_leaf_138_clk),
    .Q(\register_file[22][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16268_ (.D(_00656_),
    .CLK(clknet_leaf_138_clk),
    .Q(\register_file[22][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16269_ (.D(_00657_),
    .CLK(clknet_leaf_139_clk),
    .Q(\register_file[22][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16270_ (.D(_00658_),
    .CLK(clknet_leaf_153_clk),
    .Q(\register_file[22][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16271_ (.D(_00659_),
    .CLK(clknet_leaf_154_clk),
    .Q(\register_file[22][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16272_ (.D(_00660_),
    .CLK(clknet_leaf_155_clk),
    .Q(\register_file[22][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16273_ (.D(_00661_),
    .CLK(clknet_leaf_158_clk),
    .Q(\register_file[22][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16274_ (.D(_00662_),
    .CLK(clknet_leaf_158_clk),
    .Q(\register_file[22][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16275_ (.D(_00663_),
    .CLK(clknet_leaf_209_clk),
    .Q(\register_file[22][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16276_ (.D(_00664_),
    .CLK(clknet_leaf_208_clk),
    .Q(\register_file[22][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16277_ (.D(_00665_),
    .CLK(clknet_leaf_208_clk),
    .Q(\register_file[22][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16278_ (.D(_00666_),
    .CLK(clknet_leaf_207_clk),
    .Q(\register_file[22][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16279_ (.D(_00667_),
    .CLK(clknet_leaf_197_clk),
    .Q(\register_file[22][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16280_ (.D(_00668_),
    .CLK(clknet_leaf_191_clk),
    .Q(\register_file[22][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16281_ (.D(_00669_),
    .CLK(clknet_leaf_193_clk),
    .Q(\register_file[22][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16282_ (.D(_00670_),
    .CLK(clknet_leaf_269_clk),
    .Q(\register_file[22][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16283_ (.D(_00671_),
    .CLK(clknet_leaf_40_clk),
    .Q(\register_file[22][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16284_ (.D(_00672_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\register_file[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16285_ (.D(_00673_),
    .CLK(clknet_leaf_30_clk),
    .Q(\register_file[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16286_ (.D(_00674_),
    .CLK(clknet_leaf_27_clk),
    .Q(\register_file[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16287_ (.D(_00675_),
    .CLK(clknet_leaf_17_clk),
    .Q(\register_file[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16288_ (.D(_00676_),
    .CLK(clknet_leaf_16_clk),
    .Q(\register_file[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16289_ (.D(_00677_),
    .CLK(clknet_leaf_68_clk),
    .Q(\register_file[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16290_ (.D(_00678_),
    .CLK(clknet_leaf_68_clk),
    .Q(\register_file[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16291_ (.D(_00679_),
    .CLK(clknet_leaf_68_clk),
    .Q(\register_file[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16292_ (.D(_00680_),
    .CLK(clknet_leaf_74_clk),
    .Q(\register_file[21][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16293_ (.D(_00681_),
    .CLK(clknet_leaf_75_clk),
    .Q(\register_file[21][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16294_ (.D(_00682_),
    .CLK(clknet_leaf_80_clk),
    .Q(\register_file[21][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16295_ (.D(_00683_),
    .CLK(clknet_leaf_80_clk),
    .Q(\register_file[21][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16296_ (.D(_00684_),
    .CLK(clknet_leaf_80_clk),
    .Q(\register_file[21][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16297_ (.D(_00685_),
    .CLK(clknet_leaf_97_clk),
    .Q(\register_file[21][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16298_ (.D(_00686_),
    .CLK(clknet_leaf_97_clk),
    .Q(\register_file[21][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16299_ (.D(_00687_),
    .CLK(clknet_leaf_138_clk),
    .Q(\register_file[21][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16300_ (.D(_00688_),
    .CLK(clknet_leaf_139_clk),
    .Q(\register_file[21][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16301_ (.D(_00689_),
    .CLK(clknet_leaf_143_clk),
    .Q(\register_file[21][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16302_ (.D(_00690_),
    .CLK(clknet_leaf_145_clk),
    .Q(\register_file[21][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16303_ (.D(_00691_),
    .CLK(clknet_leaf_145_clk),
    .Q(\register_file[21][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16304_ (.D(_00692_),
    .CLK(clknet_leaf_158_clk),
    .Q(\register_file[21][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16305_ (.D(_00693_),
    .CLK(clknet_leaf_159_clk),
    .Q(\register_file[21][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16306_ (.D(_00694_),
    .CLK(clknet_leaf_158_clk),
    .Q(\register_file[21][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16307_ (.D(_00695_),
    .CLK(clknet_leaf_209_clk),
    .Q(\register_file[21][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16308_ (.D(_00696_),
    .CLK(clknet_leaf_180_clk),
    .Q(\register_file[21][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16309_ (.D(_00697_),
    .CLK(clknet_leaf_206_clk),
    .Q(\register_file[21][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16310_ (.D(_00698_),
    .CLK(clknet_leaf_182_clk),
    .Q(\register_file[21][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16311_ (.D(_00699_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\register_file[21][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16312_ (.D(_00700_),
    .CLK(clknet_leaf_194_clk),
    .Q(\register_file[21][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16313_ (.D(_00701_),
    .CLK(clknet_leaf_194_clk),
    .Q(\register_file[21][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16314_ (.D(_00702_),
    .CLK(clknet_leaf_270_clk),
    .Q(\register_file[21][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16315_ (.D(_00703_),
    .CLK(clknet_leaf_272_clk),
    .Q(\register_file[21][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16316_ (.D(_00704_),
    .CLK(clknet_leaf_278_clk),
    .Q(\register_file[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16317_ (.D(_00705_),
    .CLK(clknet_leaf_30_clk),
    .Q(\register_file[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16318_ (.D(_00706_),
    .CLK(clknet_leaf_30_clk),
    .Q(\register_file[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16319_ (.D(_00707_),
    .CLK(clknet_leaf_15_clk),
    .Q(\register_file[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16320_ (.D(_00708_),
    .CLK(clknet_leaf_19_clk),
    .Q(\register_file[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16321_ (.D(_00709_),
    .CLK(clknet_leaf_67_clk),
    .Q(\register_file[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16322_ (.D(_00710_),
    .CLK(clknet_leaf_60_clk),
    .Q(\register_file[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16323_ (.D(_00711_),
    .CLK(clknet_leaf_68_clk),
    .Q(\register_file[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16324_ (.D(_00712_),
    .CLK(clknet_leaf_73_clk),
    .Q(\register_file[20][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16325_ (.D(_00713_),
    .CLK(clknet_leaf_77_clk),
    .Q(\register_file[20][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16326_ (.D(_00714_),
    .CLK(clknet_leaf_81_clk),
    .Q(\register_file[20][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16327_ (.D(_00715_),
    .CLK(clknet_leaf_80_clk),
    .Q(\register_file[20][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16328_ (.D(_00716_),
    .CLK(clknet_leaf_79_clk),
    .Q(\register_file[20][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16329_ (.D(_00717_),
    .CLK(clknet_leaf_99_clk),
    .Q(\register_file[20][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16330_ (.D(_00718_),
    .CLK(clknet_leaf_99_clk),
    .Q(\register_file[20][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16331_ (.D(_00719_),
    .CLK(clknet_leaf_137_clk),
    .Q(\register_file[20][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16332_ (.D(_00720_),
    .CLK(clknet_leaf_141_clk),
    .Q(\register_file[20][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16333_ (.D(_00721_),
    .CLK(clknet_leaf_142_clk),
    .Q(\register_file[20][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16334_ (.D(_00722_),
    .CLK(clknet_leaf_145_clk),
    .Q(\register_file[20][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16335_ (.D(_00723_),
    .CLK(clknet_leaf_146_clk),
    .Q(\register_file[20][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16336_ (.D(_00724_),
    .CLK(clknet_leaf_162_clk),
    .Q(\register_file[20][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16337_ (.D(_00725_),
    .CLK(clknet_leaf_157_clk),
    .Q(\register_file[20][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16338_ (.D(_00726_),
    .CLK(clknet_leaf_162_clk),
    .Q(\register_file[20][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16339_ (.D(_00727_),
    .CLK(clknet_leaf_210_clk),
    .Q(\register_file[20][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16340_ (.D(_00728_),
    .CLK(clknet_leaf_180_clk),
    .Q(\register_file[20][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16341_ (.D(_00729_),
    .CLK(clknet_leaf_206_clk),
    .Q(\register_file[20][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16342_ (.D(_00730_),
    .CLK(clknet_leaf_182_clk),
    .Q(\register_file[20][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16343_ (.D(_00731_),
    .CLK(clknet_leaf_197_clk),
    .Q(\register_file[20][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16344_ (.D(_00732_),
    .CLK(clknet_leaf_195_clk),
    .Q(\register_file[20][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16345_ (.D(_00733_),
    .CLK(clknet_leaf_196_clk),
    .Q(\register_file[20][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16346_ (.D(_00734_),
    .CLK(clknet_leaf_270_clk),
    .Q(\register_file[20][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16347_ (.D(_00735_),
    .CLK(clknet_leaf_272_clk),
    .Q(\register_file[20][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16348_ (.D(_00736_),
    .CLK(clknet_leaf_281_clk),
    .Q(\register_file[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16349_ (.D(_00737_),
    .CLK(clknet_leaf_302_clk),
    .Q(\register_file[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16350_ (.D(_00738_),
    .CLK(clknet_leaf_303_clk),
    .Q(\register_file[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16351_ (.D(_00739_),
    .CLK(clknet_leaf_3_clk),
    .Q(\register_file[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16352_ (.D(_00740_),
    .CLK(clknet_leaf_3_clk),
    .Q(\register_file[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16353_ (.D(_00741_),
    .CLK(clknet_leaf_58_clk),
    .Q(\register_file[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16354_ (.D(_00742_),
    .CLK(clknet_leaf_58_clk),
    .Q(\register_file[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16355_ (.D(_00743_),
    .CLK(clknet_leaf_58_clk),
    .Q(\register_file[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16356_ (.D(_00744_),
    .CLK(clknet_leaf_74_clk),
    .Q(\register_file[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16357_ (.D(_00745_),
    .CLK(clknet_leaf_74_clk),
    .Q(\register_file[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16358_ (.D(_00746_),
    .CLK(clknet_leaf_82_clk),
    .Q(\register_file[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16359_ (.D(_00747_),
    .CLK(clknet_leaf_82_clk),
    .Q(\register_file[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16360_ (.D(_00748_),
    .CLK(clknet_leaf_82_clk),
    .Q(\register_file[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16361_ (.D(_00749_),
    .CLK(clknet_leaf_96_clk),
    .Q(\register_file[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16362_ (.D(_00750_),
    .CLK(clknet_leaf_96_clk),
    .Q(\register_file[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16363_ (.D(_00751_),
    .CLK(clknet_leaf_140_clk),
    .Q(\register_file[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16364_ (.D(_00752_),
    .CLK(clknet_leaf_140_clk),
    .Q(\register_file[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16365_ (.D(_00753_),
    .CLK(clknet_leaf_143_clk),
    .Q(\register_file[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16366_ (.D(_00754_),
    .CLK(clknet_leaf_144_clk),
    .Q(\register_file[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16367_ (.D(_00755_),
    .CLK(clknet_leaf_144_clk),
    .Q(\register_file[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16368_ (.D(_00756_),
    .CLK(clknet_leaf_161_clk),
    .Q(\register_file[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16369_ (.D(_00757_),
    .CLK(clknet_leaf_160_clk),
    .Q(\register_file[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16370_ (.D(_00758_),
    .CLK(clknet_leaf_159_clk),
    .Q(\register_file[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16371_ (.D(_00759_),
    .CLK(clknet_leaf_211_clk),
    .Q(\register_file[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16372_ (.D(_00760_),
    .CLK(clknet_leaf_209_clk),
    .Q(\register_file[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16373_ (.D(_00761_),
    .CLK(clknet_leaf_222_clk),
    .Q(\register_file[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16374_ (.D(_00762_),
    .CLK(clknet_leaf_223_clk),
    .Q(\register_file[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16375_ (.D(_00763_),
    .CLK(clknet_leaf_202_clk),
    .Q(\register_file[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16376_ (.D(_00764_),
    .CLK(clknet_leaf_240_clk),
    .Q(\register_file[1][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16377_ (.D(_00765_),
    .CLK(clknet_leaf_202_clk),
    .Q(\register_file[1][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16378_ (.D(_00766_),
    .CLK(clknet_leaf_255_clk),
    .Q(\register_file[1][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16379_ (.D(_00767_),
    .CLK(clknet_leaf_284_clk),
    .Q(\register_file[1][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16380_ (.D(_00768_),
    .CLK(clknet_leaf_278_clk),
    .Q(\register_file[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16381_ (.D(_00769_),
    .CLK(clknet_leaf_29_clk),
    .Q(\register_file[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16382_ (.D(_00770_),
    .CLK(clknet_leaf_29_clk),
    .Q(\register_file[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16383_ (.D(_00771_),
    .CLK(clknet_leaf_15_clk),
    .Q(\register_file[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16384_ (.D(_00772_),
    .CLK(clknet_leaf_17_clk),
    .Q(\register_file[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16385_ (.D(_00773_),
    .CLK(clknet_leaf_59_clk),
    .Q(\register_file[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16386_ (.D(_00774_),
    .CLK(clknet_leaf_60_clk),
    .Q(\register_file[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16387_ (.D(_00775_),
    .CLK(clknet_leaf_60_clk),
    .Q(\register_file[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16388_ (.D(_00776_),
    .CLK(clknet_leaf_75_clk),
    .Q(\register_file[18][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16389_ (.D(_00777_),
    .CLK(clknet_leaf_74_clk),
    .Q(\register_file[18][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16390_ (.D(_00778_),
    .CLK(clknet_leaf_82_clk),
    .Q(\register_file[18][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16391_ (.D(_00779_),
    .CLK(clknet_leaf_82_clk),
    .Q(\register_file[18][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16392_ (.D(_00780_),
    .CLK(clknet_leaf_82_clk),
    .Q(\register_file[18][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16393_ (.D(_00781_),
    .CLK(clknet_leaf_97_clk),
    .Q(\register_file[18][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16394_ (.D(_00782_),
    .CLK(clknet_leaf_97_clk),
    .Q(\register_file[18][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16395_ (.D(_00783_),
    .CLK(clknet_leaf_139_clk),
    .Q(\register_file[18][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16396_ (.D(_00784_),
    .CLK(clknet_leaf_140_clk),
    .Q(\register_file[18][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16397_ (.D(_00785_),
    .CLK(clknet_leaf_142_clk),
    .Q(\register_file[18][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16398_ (.D(_00786_),
    .CLK(clknet_leaf_144_clk),
    .Q(\register_file[18][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16399_ (.D(_00787_),
    .CLK(clknet_leaf_144_clk),
    .Q(\register_file[18][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16400_ (.D(_00788_),
    .CLK(clknet_leaf_160_clk),
    .Q(\register_file[18][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16401_ (.D(_00789_),
    .CLK(clknet_leaf_160_clk),
    .Q(\register_file[18][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16402_ (.D(_00790_),
    .CLK(clknet_leaf_159_clk),
    .Q(\register_file[18][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16403_ (.D(_00791_),
    .CLK(clknet_leaf_168_clk),
    .Q(\register_file[18][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16404_ (.D(_00792_),
    .CLK(clknet_leaf_173_clk),
    .Q(\register_file[18][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16405_ (.D(_00793_),
    .CLK(clknet_leaf_213_clk),
    .Q(\register_file[18][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16406_ (.D(_00794_),
    .CLK(clknet_leaf_214_clk),
    .Q(\register_file[18][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16407_ (.D(_00795_),
    .CLK(clknet_leaf_201_clk),
    .Q(\register_file[18][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16408_ (.D(_00796_),
    .CLK(clknet_leaf_195_clk),
    .Q(\register_file[18][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16409_ (.D(_00797_),
    .CLK(clknet_leaf_263_clk),
    .Q(\register_file[18][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16410_ (.D(_00798_),
    .CLK(clknet_leaf_272_clk),
    .Q(\register_file[18][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16411_ (.D(_00799_),
    .CLK(clknet_leaf_277_clk),
    .Q(\register_file[18][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16412_ (.D(_00800_),
    .CLK(clknet_leaf_277_clk),
    .Q(\register_file[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16413_ (.D(_00801_),
    .CLK(clknet_leaf_28_clk),
    .Q(\register_file[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16414_ (.D(_00802_),
    .CLK(clknet_leaf_27_clk),
    .Q(\register_file[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16415_ (.D(_00803_),
    .CLK(clknet_leaf_15_clk),
    .Q(\register_file[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16416_ (.D(_00804_),
    .CLK(clknet_leaf_15_clk),
    .Q(\register_file[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16417_ (.D(_00805_),
    .CLK(clknet_leaf_59_clk),
    .Q(\register_file[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16418_ (.D(_00806_),
    .CLK(clknet_leaf_59_clk),
    .Q(\register_file[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16419_ (.D(_00807_),
    .CLK(clknet_leaf_59_clk),
    .Q(\register_file[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16420_ (.D(_00808_),
    .CLK(clknet_leaf_73_clk),
    .Q(\register_file[17][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16421_ (.D(_00809_),
    .CLK(clknet_leaf_73_clk),
    .Q(\register_file[17][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16422_ (.D(_00810_),
    .CLK(clknet_leaf_83_clk),
    .Q(\register_file[17][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16423_ (.D(_00811_),
    .CLK(clknet_leaf_81_clk),
    .Q(\register_file[17][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16424_ (.D(_00812_),
    .CLK(clknet_leaf_83_clk),
    .Q(\register_file[17][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16425_ (.D(_00813_),
    .CLK(clknet_leaf_99_clk),
    .Q(\register_file[17][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16426_ (.D(_00814_),
    .CLK(clknet_leaf_98_clk),
    .Q(\register_file[17][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16427_ (.D(_00815_),
    .CLK(clknet_leaf_141_clk),
    .Q(\register_file[17][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16428_ (.D(_00816_),
    .CLK(clknet_leaf_140_clk),
    .Q(\register_file[17][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16429_ (.D(_00817_),
    .CLK(clknet_leaf_142_clk),
    .Q(\register_file[17][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16430_ (.D(_00818_),
    .CLK(clknet_leaf_147_clk),
    .Q(\register_file[17][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16431_ (.D(_00819_),
    .CLK(clknet_leaf_144_clk),
    .Q(\register_file[17][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16432_ (.D(_00820_),
    .CLK(clknet_leaf_161_clk),
    .Q(\register_file[17][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16433_ (.D(_00821_),
    .CLK(clknet_leaf_162_clk),
    .Q(\register_file[17][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16434_ (.D(_00822_),
    .CLK(clknet_leaf_165_clk),
    .Q(\register_file[17][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16435_ (.D(_00823_),
    .CLK(clknet_leaf_167_clk),
    .Q(\register_file[17][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16436_ (.D(_00824_),
    .CLK(clknet_leaf_167_clk),
    .Q(\register_file[17][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16437_ (.D(_00825_),
    .CLK(clknet_leaf_205_clk),
    .Q(\register_file[17][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16438_ (.D(_00826_),
    .CLK(clknet_leaf_204_clk),
    .Q(\register_file[17][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16439_ (.D(_00827_),
    .CLK(clknet_leaf_204_clk),
    .Q(\register_file[17][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16440_ (.D(_00828_),
    .CLK(clknet_leaf_204_clk),
    .Q(\register_file[17][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16441_ (.D(_00829_),
    .CLK(clknet_leaf_201_clk),
    .Q(\register_file[17][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16442_ (.D(_00830_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\register_file[17][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16443_ (.D(_00831_),
    .CLK(clknet_leaf_274_clk),
    .Q(\register_file[17][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16444_ (.D(_00832_),
    .CLK(clknet_leaf_286_clk),
    .Q(\register_file[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16445_ (.D(_00833_),
    .CLK(clknet_leaf_304_clk),
    .Q(\register_file[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16446_ (.D(_00834_),
    .CLK(clknet_leaf_304_clk),
    .Q(\register_file[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16447_ (.D(_00835_),
    .CLK(clknet_leaf_2_clk),
    .Q(\register_file[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16448_ (.D(_00836_),
    .CLK(clknet_leaf_2_clk),
    .Q(\register_file[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16449_ (.D(_00837_),
    .CLK(clknet_leaf_54_clk),
    .Q(\register_file[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16450_ (.D(_00838_),
    .CLK(clknet_leaf_52_clk),
    .Q(\register_file[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16451_ (.D(_00839_),
    .CLK(clknet_leaf_56_clk),
    .Q(\register_file[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16452_ (.D(_00840_),
    .CLK(clknet_leaf_67_clk),
    .Q(\register_file[16][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16453_ (.D(_00841_),
    .CLK(clknet_leaf_67_clk),
    .Q(\register_file[16][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16454_ (.D(_00842_),
    .CLK(clknet_leaf_86_clk),
    .Q(\register_file[16][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16455_ (.D(_00843_),
    .CLK(clknet_leaf_64_clk),
    .Q(\register_file[16][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16456_ (.D(_00844_),
    .CLK(clknet_leaf_86_clk),
    .Q(\register_file[16][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16457_ (.D(_00845_),
    .CLK(clknet_leaf_104_clk),
    .Q(\register_file[16][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16458_ (.D(_00846_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\register_file[16][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16459_ (.D(_00847_),
    .CLK(clknet_leaf_130_clk),
    .Q(\register_file[16][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16460_ (.D(_00848_),
    .CLK(clknet_leaf_131_clk),
    .Q(\register_file[16][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16461_ (.D(_00849_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\register_file[16][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16462_ (.D(_00850_),
    .CLK(clknet_leaf_129_clk),
    .Q(\register_file[16][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16463_ (.D(_00851_),
    .CLK(clknet_leaf_148_clk),
    .Q(\register_file[16][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16464_ (.D(_00852_),
    .CLK(clknet_leaf_166_clk),
    .Q(\register_file[16][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16465_ (.D(_00853_),
    .CLK(clknet_leaf_164_clk),
    .Q(\register_file[16][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16466_ (.D(_00854_),
    .CLK(clknet_leaf_166_clk),
    .Q(\register_file[16][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16467_ (.D(_00855_),
    .CLK(clknet_leaf_167_clk),
    .Q(\register_file[16][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16468_ (.D(_00856_),
    .CLK(clknet_leaf_167_clk),
    .Q(\register_file[16][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16469_ (.D(_00857_),
    .CLK(clknet_leaf_215_clk),
    .Q(\register_file[16][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16470_ (.D(_00858_),
    .CLK(clknet_leaf_216_clk),
    .Q(\register_file[16][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16471_ (.D(_00859_),
    .CLK(clknet_leaf_215_clk),
    .Q(\register_file[16][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16472_ (.D(_00860_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\register_file[16][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16473_ (.D(_00861_),
    .CLK(clknet_leaf_202_clk),
    .Q(\register_file[16][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16474_ (.D(_00862_),
    .CLK(clknet_leaf_253_clk),
    .Q(\register_file[16][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16475_ (.D(_00863_),
    .CLK(clknet_leaf_285_clk),
    .Q(\register_file[16][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16476_ (.D(_00864_),
    .CLK(clknet_leaf_282_clk),
    .Q(\register_file[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16477_ (.D(_00865_),
    .CLK(clknet_leaf_301_clk),
    .Q(\register_file[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16478_ (.D(_00866_),
    .CLK(clknet_leaf_305_clk),
    .Q(\register_file[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16479_ (.D(_00867_),
    .CLK(clknet_leaf_6_clk),
    .Q(\register_file[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16480_ (.D(_00868_),
    .CLK(clknet_leaf_6_clk),
    .Q(\register_file[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16481_ (.D(_00869_),
    .CLK(clknet_leaf_22_clk),
    .Q(\register_file[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16482_ (.D(_00870_),
    .CLK(clknet_leaf_53_clk),
    .Q(\register_file[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16483_ (.D(_00871_),
    .CLK(clknet_leaf_52_clk),
    .Q(\register_file[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16484_ (.D(_00872_),
    .CLK(clknet_leaf_57_clk),
    .Q(\register_file[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16485_ (.D(_00873_),
    .CLK(clknet_leaf_61_clk),
    .Q(\register_file[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16486_ (.D(_00874_),
    .CLK(clknet_leaf_48_clk),
    .Q(\register_file[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16487_ (.D(_00875_),
    .CLK(clknet_leaf_48_clk),
    .Q(\register_file[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16488_ (.D(_00876_),
    .CLK(clknet_leaf_48_clk),
    .Q(\register_file[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16489_ (.D(_00877_),
    .CLK(clknet_leaf_110_clk),
    .Q(\register_file[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16490_ (.D(_00878_),
    .CLK(clknet_leaf_114_clk),
    .Q(\register_file[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16491_ (.D(_00879_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\register_file[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16492_ (.D(_00880_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\register_file[15][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16493_ (.D(_00881_),
    .CLK(clknet_leaf_125_clk),
    .Q(\register_file[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16494_ (.D(_00882_),
    .CLK(clknet_leaf_188_clk),
    .Q(\register_file[15][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16495_ (.D(_00883_),
    .CLK(clknet_leaf_188_clk),
    .Q(\register_file[15][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16496_ (.D(_00884_),
    .CLK(clknet_leaf_174_clk),
    .Q(\register_file[15][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16497_ (.D(_00885_),
    .CLK(clknet_leaf_175_clk),
    .Q(\register_file[15][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16498_ (.D(_00886_),
    .CLK(clknet_leaf_175_clk),
    .Q(\register_file[15][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16499_ (.D(_00887_),
    .CLK(clknet_leaf_174_clk),
    .Q(\register_file[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16500_ (.D(_00888_),
    .CLK(clknet_leaf_174_clk),
    .Q(\register_file[15][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16501_ (.D(_00889_),
    .CLK(clknet_leaf_225_clk),
    .Q(\register_file[15][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16502_ (.D(_00890_),
    .CLK(clknet_leaf_225_clk),
    .Q(\register_file[15][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16503_ (.D(_00891_),
    .CLK(clknet_leaf_222_clk),
    .Q(\register_file[15][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16504_ (.D(_00892_),
    .CLK(clknet_leaf_242_clk),
    .Q(\register_file[15][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16505_ (.D(_00893_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\register_file[15][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16506_ (.D(_00894_),
    .CLK(clknet_leaf_254_clk),
    .Q(\register_file[15][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16507_ (.D(_00895_),
    .CLK(clknet_leaf_286_clk),
    .Q(\register_file[15][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16508_ (.D(_00896_),
    .CLK(clknet_leaf_287_clk),
    .Q(\register_file[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16509_ (.D(_00897_),
    .CLK(clknet_leaf_300_clk),
    .Q(\register_file[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16510_ (.D(_00898_),
    .CLK(clknet_leaf_305_clk),
    .Q(\register_file[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16511_ (.D(_00899_),
    .CLK(clknet_leaf_2_clk),
    .Q(\register_file[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16512_ (.D(_00900_),
    .CLK(clknet_leaf_1_clk),
    .Q(\register_file[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16513_ (.D(_00901_),
    .CLK(clknet_leaf_22_clk),
    .Q(\register_file[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16514_ (.D(_00902_),
    .CLK(clknet_leaf_20_clk),
    .Q(\register_file[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16515_ (.D(_00903_),
    .CLK(clknet_leaf_22_clk),
    .Q(\register_file[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16516_ (.D(_00904_),
    .CLK(clknet_leaf_59_clk),
    .Q(\register_file[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16517_ (.D(_00905_),
    .CLK(clknet_leaf_59_clk),
    .Q(\register_file[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16518_ (.D(_00906_),
    .CLK(clknet_leaf_48_clk),
    .Q(\register_file[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16519_ (.D(_00907_),
    .CLK(clknet_leaf_48_clk),
    .Q(\register_file[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16520_ (.D(_00908_),
    .CLK(clknet_leaf_46_clk),
    .Q(\register_file[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16521_ (.D(_00909_),
    .CLK(clknet_leaf_110_clk),
    .Q(\register_file[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16522_ (.D(_00910_),
    .CLK(clknet_leaf_110_clk),
    .Q(\register_file[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16523_ (.D(_00911_),
    .CLK(clknet_leaf_124_clk),
    .Q(\register_file[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16524_ (.D(_00912_),
    .CLK(clknet_leaf_123_clk),
    .Q(\register_file[14][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16525_ (.D(_00913_),
    .CLK(clknet_leaf_125_clk),
    .Q(\register_file[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16526_ (.D(_00914_),
    .CLK(clknet_leaf_125_clk),
    .Q(\register_file[14][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16527_ (.D(_00915_),
    .CLK(clknet_leaf_126_clk),
    .Q(\register_file[14][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16528_ (.D(_00916_),
    .CLK(clknet_leaf_173_clk),
    .Q(\register_file[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16529_ (.D(_00917_),
    .CLK(clknet_leaf_172_clk),
    .Q(\register_file[14][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16530_ (.D(_00918_),
    .CLK(clknet_leaf_175_clk),
    .Q(\register_file[14][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16531_ (.D(_00919_),
    .CLK(clknet_leaf_174_clk),
    .Q(\register_file[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16532_ (.D(_00920_),
    .CLK(clknet_leaf_174_clk),
    .Q(\register_file[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16533_ (.D(_00921_),
    .CLK(clknet_leaf_225_clk),
    .Q(\register_file[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16534_ (.D(_00922_),
    .CLK(clknet_leaf_226_clk),
    .Q(\register_file[14][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16535_ (.D(_00923_),
    .CLK(clknet_leaf_226_clk),
    .Q(\register_file[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16536_ (.D(_00924_),
    .CLK(clknet_leaf_241_clk),
    .Q(\register_file[14][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16537_ (.D(_00925_),
    .CLK(clknet_leaf_241_clk),
    .Q(\register_file[14][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16538_ (.D(_00926_),
    .CLK(clknet_leaf_254_clk),
    .Q(\register_file[14][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16539_ (.D(_00927_),
    .CLK(clknet_leaf_287_clk),
    .Q(\register_file[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16540_ (.D(_00928_),
    .CLK(clknet_leaf_282_clk),
    .Q(\register_file[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16541_ (.D(_00929_),
    .CLK(clknet_leaf_301_clk),
    .Q(\register_file[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16542_ (.D(_00930_),
    .CLK(clknet_leaf_302_clk),
    .Q(\register_file[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16543_ (.D(_00931_),
    .CLK(clknet_leaf_4_clk),
    .Q(\register_file[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16544_ (.D(_00932_),
    .CLK(clknet_leaf_5_clk),
    .Q(\register_file[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16545_ (.D(_00933_),
    .CLK(clknet_leaf_18_clk),
    .Q(\register_file[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16546_ (.D(_00934_),
    .CLK(clknet_leaf_19_clk),
    .Q(\register_file[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16547_ (.D(_00935_),
    .CLK(clknet_leaf_18_clk),
    .Q(\register_file[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16548_ (.D(_00936_),
    .CLK(clknet_leaf_69_clk),
    .Q(\register_file[29][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16549_ (.D(_00937_),
    .CLK(clknet_leaf_65_clk),
    .Q(\register_file[29][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16550_ (.D(_00938_),
    .CLK(clknet_leaf_85_clk),
    .Q(\register_file[29][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16551_ (.D(_00939_),
    .CLK(clknet_leaf_85_clk),
    .Q(\register_file[29][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16552_ (.D(_00940_),
    .CLK(clknet_leaf_85_clk),
    .Q(\register_file[29][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16553_ (.D(_00941_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\register_file[29][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16554_ (.D(_00942_),
    .CLK(clknet_leaf_105_clk),
    .Q(\register_file[29][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16555_ (.D(_00943_),
    .CLK(clknet_leaf_134_clk),
    .Q(\register_file[29][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16556_ (.D(_00944_),
    .CLK(clknet_leaf_130_clk),
    .Q(\register_file[29][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16557_ (.D(_00945_),
    .CLK(clknet_leaf_129_clk),
    .Q(\register_file[29][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16558_ (.D(_00946_),
    .CLK(clknet_leaf_150_clk),
    .Q(\register_file[29][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16559_ (.D(_00947_),
    .CLK(clknet_leaf_150_clk),
    .Q(\register_file[29][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16560_ (.D(_00948_),
    .CLK(clknet_leaf_164_clk),
    .Q(\register_file[29][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16561_ (.D(_00949_),
    .CLK(clknet_leaf_165_clk),
    .Q(\register_file[29][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16562_ (.D(_00950_),
    .CLK(clknet_leaf_180_clk),
    .Q(\register_file[29][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16563_ (.D(_00951_),
    .CLK(clknet_leaf_179_clk),
    .Q(\register_file[29][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16564_ (.D(_00952_),
    .CLK(clknet_leaf_210_clk),
    .Q(\register_file[29][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16565_ (.D(_00953_),
    .CLK(clknet_leaf_215_clk),
    .Q(\register_file[29][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16566_ (.D(_00954_),
    .CLK(clknet_leaf_215_clk),
    .Q(\register_file[29][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16567_ (.D(_00955_),
    .CLK(clknet_leaf_215_clk),
    .Q(\register_file[29][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16568_ (.D(_00956_),
    .CLK(clknet_leaf_262_clk),
    .Q(\register_file[29][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16569_ (.D(_00957_),
    .CLK(clknet_leaf_263_clk),
    .Q(\register_file[29][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16570_ (.D(_00958_),
    .CLK(clknet_leaf_253_clk),
    .Q(\register_file[29][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16571_ (.D(_00959_),
    .CLK(clknet_leaf_285_clk),
    .Q(\register_file[29][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16572_ (.D(_00960_),
    .CLK(clknet_leaf_286_clk),
    .Q(\register_file[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16573_ (.D(_00961_),
    .CLK(clknet_leaf_304_clk),
    .Q(\register_file[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16574_ (.D(_00962_),
    .CLK(clknet_leaf_305_clk),
    .Q(\register_file[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16575_ (.D(_00963_),
    .CLK(clknet_leaf_5_clk),
    .Q(\register_file[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16576_ (.D(_00964_),
    .CLK(clknet_leaf_5_clk),
    .Q(\register_file[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16577_ (.D(_00965_),
    .CLK(clknet_leaf_14_clk),
    .Q(\register_file[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16578_ (.D(_00966_),
    .CLK(clknet_leaf_14_clk),
    .Q(\register_file[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16579_ (.D(_00967_),
    .CLK(clknet_leaf_13_clk),
    .Q(\register_file[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16580_ (.D(_00968_),
    .CLK(clknet_leaf_57_clk),
    .Q(\register_file[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16581_ (.D(_00969_),
    .CLK(clknet_leaf_57_clk),
    .Q(\register_file[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16582_ (.D(_00970_),
    .CLK(clknet_leaf_49_clk),
    .Q(\register_file[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16583_ (.D(_00971_),
    .CLK(clknet_leaf_49_clk),
    .Q(\register_file[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16584_ (.D(_00972_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\register_file[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16585_ (.D(_00973_),
    .CLK(clknet_leaf_114_clk),
    .Q(\register_file[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16586_ (.D(_00974_),
    .CLK(clknet_leaf_115_clk),
    .Q(\register_file[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16587_ (.D(_00975_),
    .CLK(clknet_leaf_115_clk),
    .Q(\register_file[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16588_ (.D(_00976_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\register_file[9][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16589_ (.D(_00977_),
    .CLK(clknet_leaf_117_clk),
    .Q(\register_file[9][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16590_ (.D(_00978_),
    .CLK(clknet_leaf_188_clk),
    .Q(\register_file[9][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16591_ (.D(_00979_),
    .CLK(clknet_leaf_189_clk),
    .Q(\register_file[9][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16592_ (.D(_00980_),
    .CLK(clknet_leaf_176_clk),
    .Q(\register_file[9][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16593_ (.D(_00981_),
    .CLK(clknet_leaf_178_clk),
    .Q(\register_file[9][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16594_ (.D(_00982_),
    .CLK(clknet_leaf_176_clk),
    .Q(\register_file[9][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16595_ (.D(_00983_),
    .CLK(clknet_leaf_214_clk),
    .Q(\register_file[9][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16596_ (.D(_00984_),
    .CLK(clknet_leaf_214_clk),
    .Q(\register_file[9][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16597_ (.D(_00985_),
    .CLK(clknet_leaf_217_clk),
    .Q(\register_file[9][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16598_ (.D(_00986_),
    .CLK(clknet_leaf_224_clk),
    .Q(\register_file[9][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16599_ (.D(_00987_),
    .CLK(clknet_leaf_223_clk),
    .Q(\register_file[9][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16600_ (.D(_00988_),
    .CLK(clknet_leaf_257_clk),
    .Q(\register_file[9][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16601_ (.D(_00989_),
    .CLK(clknet_leaf_257_clk),
    .Q(\register_file[9][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16602_ (.D(_00990_),
    .CLK(clknet_leaf_253_clk),
    .Q(\register_file[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16603_ (.D(_00991_),
    .CLK(clknet_leaf_284_clk),
    .Q(\register_file[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1 (.I(addrD[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(addrD[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(addrD[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(addrD[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(addrD[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(addrS[0]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(addrS[1]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(addrS[2]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(addrS[3]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(addrS[4]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(new_value[0]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(new_value[10]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(new_value[11]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(new_value[12]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(new_value[13]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(new_value[14]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(new_value[15]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(new_value[16]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(new_value[17]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(new_value[18]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(new_value[19]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(new_value[1]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(new_value[20]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(new_value[21]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(new_value[22]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(new_value[23]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(new_value[24]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(new_value[25]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(new_value[26]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(new_value[27]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(new_value[28]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(new_value[29]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(new_value[2]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(new_value[30]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(new_value[31]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(new_value[3]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(new_value[4]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(new_value[5]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(new_value[6]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(new_value[7]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(new_value[8]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(new_value[9]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(we),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output44 (.I(net44),
    .Z(rD[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output45 (.I(net45),
    .Z(rD[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output46 (.I(net46),
    .Z(rD[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output47 (.I(net47),
    .Z(rD[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output48 (.I(net48),
    .Z(rD[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output49 (.I(net49),
    .Z(rD[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output50 (.I(net50),
    .Z(rD[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output51 (.I(net51),
    .Z(rD[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output52 (.I(net52),
    .Z(rD[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output53 (.I(net53),
    .Z(rD[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output54 (.I(net54),
    .Z(rD[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output55 (.I(net55),
    .Z(rD[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output56 (.I(net56),
    .Z(rD[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output57 (.I(net57),
    .Z(rD[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output58 (.I(net58),
    .Z(rD[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output59 (.I(net59),
    .Z(rD[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output60 (.I(net60),
    .Z(rD[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output61 (.I(net61),
    .Z(rD[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output62 (.I(net62),
    .Z(rD[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output63 (.I(net63),
    .Z(rD[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output64 (.I(net64),
    .Z(rD[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output65 (.I(net65),
    .Z(rD[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output66 (.I(net66),
    .Z(rD[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output67 (.I(net67),
    .Z(rD[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output68 (.I(net68),
    .Z(rD[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output69 (.I(net69),
    .Z(rD[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output70 (.I(net70),
    .Z(rD[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output71 (.I(net71),
    .Z(rD[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output72 (.I(net72),
    .Z(rD[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output73 (.I(net73),
    .Z(rD[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output74 (.I(net74),
    .Z(rD[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output75 (.I(net75),
    .Z(rD[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output76 (.I(net76),
    .Z(rS[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output77 (.I(net77),
    .Z(rS[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output78 (.I(net78),
    .Z(rS[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output79 (.I(net79),
    .Z(rS[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output80 (.I(net80),
    .Z(rS[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output81 (.I(net81),
    .Z(rS[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output82 (.I(net82),
    .Z(rS[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output83 (.I(net83),
    .Z(rS[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output84 (.I(net84),
    .Z(rS[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output85 (.I(net85),
    .Z(rS[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output86 (.I(net86),
    .Z(rS[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output87 (.I(net87),
    .Z(rS[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output88 (.I(net88),
    .Z(rS[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output89 (.I(net89),
    .Z(rS[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output90 (.I(net90),
    .Z(rS[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output91 (.I(net91),
    .Z(rS[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output92 (.I(net92),
    .Z(rS[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output93 (.I(net93),
    .Z(rS[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output94 (.I(net94),
    .Z(rS[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output95 (.I(net95),
    .Z(rS[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output96 (.I(net96),
    .Z(rS[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output97 (.I(net97),
    .Z(rS[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output98 (.I(net98),
    .Z(rS[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output99 (.I(net99),
    .Z(rS[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output100 (.I(net100),
    .Z(rS[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output101 (.I(net101),
    .Z(rS[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output102 (.I(net102),
    .Z(rS[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output103 (.I(net103),
    .Z(rS[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output104 (.I(net104),
    .Z(rS[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output105 (.I(net105),
    .Z(rS[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output106 (.I(net106),
    .Z(rS[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output107 (.I(net107),
    .Z(rS[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_111_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_122_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_123_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_124_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_129_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_130_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_131_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_132_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_134_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_137_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_140_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_141_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_143_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_145_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_146_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_147_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_148_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_151_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_151_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_153_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_154_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_155_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_155_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_156_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_157_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_158_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_158_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_159_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_159_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_160_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_160_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_161_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_161_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_162_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_164_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_164_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_165_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_166_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_167_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_168_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_168_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_169_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_169_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_170_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_170_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_171_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_171_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_172_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_172_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_173_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_174_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_175_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_176_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_176_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_177_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_178_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_179_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_179_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_180_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_180_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_181_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_182_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_182_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_183_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_183_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_185_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_185_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_186_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_187_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_187_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_188_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_188_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_189_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_189_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_190_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_191_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_192_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_192_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_193_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_194_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_194_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_195_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_195_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_196_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_196_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_197_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_199_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_199_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_201_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_201_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_202_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_202_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_203_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_203_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_204_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_204_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_205_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_205_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_206_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_206_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_207_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_207_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_208_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_208_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_209_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_210_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_210_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_211_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_212_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_212_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_213_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_214_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_215_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_216_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_217_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_217_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_218_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_218_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_219_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_219_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_220_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_220_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_221_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_222_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_222_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_223_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_223_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_224_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_225_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_225_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_226_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_228_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_228_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_229_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_230_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_231_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_233_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_233_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_234_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_234_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_235_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_235_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_237_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_237_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_238_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_238_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_239_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_239_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_240_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_240_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_241_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_242_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_242_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_243_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_244_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_245_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_245_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_246_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_246_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_247_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_247_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_248_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_248_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_249_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_249_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_250_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_250_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_251_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_251_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_252_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_252_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_253_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_254_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_254_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_255_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_255_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_256_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_256_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_257_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_257_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_259_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_259_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_260_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_260_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_261_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_261_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_262_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_262_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_263_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_263_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_264_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_264_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_265_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_265_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_267_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_267_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_269_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_269_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_270_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_270_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_271_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_271_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_272_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_272_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_274_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_274_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_275_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_275_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_276_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_276_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_277_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_277_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_278_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_278_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_279_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_279_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_280_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_280_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_281_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_281_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_282_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_282_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_283_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_283_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_284_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_284_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_285_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_285_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_286_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_286_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_287_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_287_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_288_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_288_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_289_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_289_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_291_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_291_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_292_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_292_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_293_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_293_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_295_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_295_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_296_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_296_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_297_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_297_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_298_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_298_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_299_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_299_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_300_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_300_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_301_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_301_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_302_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_302_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_303_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_303_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_304_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_304_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_305_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_305_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_306_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_306_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_307_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_307_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_309_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_309_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_310_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_310_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_313_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_314_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_0__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_1__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_2__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_3__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_4__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_5__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_6__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_7__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_8__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_9__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_10__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_11__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_12__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_13__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_14__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_15__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_16__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_17__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_18__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_19__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_20__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_21__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_22__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_23__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_24__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_25__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_26__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_27__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_28__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_29__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_30__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_31__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16096__D (.I(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16173__D (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16200__D (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16297__D (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13558__I (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13508__I (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13496__I (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13472__I (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14013__I (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13640__I (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13586__I (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13534__I (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13473__I (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14969__I (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14547__I (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14120__I (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13682__I (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13474__I (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13475__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13835__I (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13788__I (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13645__I (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13537__I (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13478__I (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15458__I (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14034__I (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13657__I (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13479__I (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__I (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13948__A1 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13860__A1 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13770__A1 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13684__A1 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13480__A1 (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13664__I (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13483__I (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15552__I (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13905__I (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13593__I (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13541__I (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13484__I (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14465__I (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14037__I (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13676__A1 (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13485__I (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__I (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13950__A2 (.I(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13862__A2 (.I(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13772__A2 (.I(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13686__A2 (.I(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13486__A2 (.I(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14741__I (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13488__I (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15479__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14319__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13973__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13773__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13489__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15584__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15330__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13490__I (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13687__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13491__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A3 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__B (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15429__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13598__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13547__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13493__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14722__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14300__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13864__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13630__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13494__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13775__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13688__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13495__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15440__I (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14469__I (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14041__I (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13498__I (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__I (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13954__A1 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13866__A1 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13776__A1 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13689__A1 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13499__A1 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15291__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13625__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13530__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13501__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13503__A1 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A3 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A3 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A2 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13637__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13571__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13524__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13512__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13503__A2 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13505__I (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__B (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__B (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__B (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13955__B (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13867__B (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13777__B (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13690__B (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13506__B (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13869__I (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13676__A2 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13510__I (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A1 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A1 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13779__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13692__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13511__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15460__I (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13611__I (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13562__I (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13514__I (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__I (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14811__I (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14389__I (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13958__I (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13515__I (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A3 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13872__A2 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13781__A2 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13694__A2 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13520__A2 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A2 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15317__I (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14897__I (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14475__I (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14048__I (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13518__I (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13959__A1 (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13871__A1 (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13780__A1 (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13693__A1 (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13519__A1 (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15311__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14891__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13961__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13522__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13873__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13782__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13695__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13523__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14816__I (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14394__I (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13963__I (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13525__I (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A3 (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13875__A2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13784__A2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13698__A2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13529__A2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__A2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15528__I (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15106__I (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14684__I (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13696__I (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13527__I (.I(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13528__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14155__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13652__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13579__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13531__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13785__A3 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13699__A3 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13532__A3 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A2 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A2 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15389__I (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14483__I (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14056__I (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13535__I (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__I (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13968__A1 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13880__A1 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13787__A1 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13701__A1 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13536__A1 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15304__I (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14884__I (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14462__I (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13538__I (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__I (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13702__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13539__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A2 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A2 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15307__I (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14887__I (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13971__I (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13542__I (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__I (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13883__A2 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13792__A2 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13704__A2 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13543__A2 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A2 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15412__I (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14720__I (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13705__I (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13596__I (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13545__I (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15564__A2 (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15309__A2 (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13546__A2 (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A2 (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15565__I (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15143__I (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14232__I (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13794__I (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13548__I (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13707__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13549__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15234__I (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14814__I (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14392__I (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13551__I (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__I (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13796__A1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13708__A1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13552__A1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__A1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15610__I (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15188__I (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14043__I (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13604__I (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13554__I (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15249__I (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14829__I (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14407__I (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13977__I (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13555__I (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13889__B (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13797__B (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13709__B (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13556__B (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__B (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15262__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14842__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14420__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13559__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15570__I (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15148__I (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14727__I (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14305__I (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13560__I (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13711__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13561__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15231__I (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14327__I (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13892__I (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13563__I (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__I (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13803__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13713__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13567__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14750__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14328__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13893__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13565__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__I (.I(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13712__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13566__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A2 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15086__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14664__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14241__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13804__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13569__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13714__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13570__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15453__I (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14178__I (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13806__I (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13572__I (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__I (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15510__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15088__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13738__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13573__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13716__A2 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13578__A2 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A3 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A2 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__A2 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14667__I (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14244__I (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13808__I (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13576__I (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__I (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13715__A1 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13577__A1 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A2 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A2 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15577__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15155__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14734__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13717__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13580__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13581__A3 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A3 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A3 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A3 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A3 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13585__A2 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15260__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14840__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13678__A2 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13584__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13901__A3 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13813__A3 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13720__A3 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13585__A3 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__A2 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13681__A1 (.I(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15325__I (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14905__I (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13991__I (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13587__I (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__I (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13902__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13814__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13721__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15008__I (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14586__I (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14161__I (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13722__I (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13590__I (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13591__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15244__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14824__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14402__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13594__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13817__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13725__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13595__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13818__A2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13726__A2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13597__A2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__A2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15499__I (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15077__I (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14655__I (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13727__I (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13599__I (.I(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13600__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15508__I (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14593__I (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14169__I (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13729__I (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13602__I (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13603__A1 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A1 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A1 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A1 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A1 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14768__I (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14346__I (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13913__I (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13605__I (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__I (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13821__B (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13731__B (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13606__B (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__B (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__B (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15019__I (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14597__I (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14173__I (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13733__I (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13609__I (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13610__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15591__I (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15169__I (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14749__I (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13824__I (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13612__I (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13736__A2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13616__A2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15592__I (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15170__I (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14262__I (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13825__I (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13614__I (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13735__A1 (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13615__A1 (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A1 (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A1 (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A1 (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15436__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15015__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14087__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13618__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14004__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13919__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13828__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13737__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13619__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13624__A2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15511__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15089__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14516__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14089__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13622__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14005__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13920__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13829__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13739__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13623__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14871__I (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14449__I (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14021__I (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13876__I (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13626__I (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15361__I (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14941__I (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14519__I (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14092__I (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13627__I (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__A3 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13922__A3 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13831__A3 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13741__A3 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13628__A3 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13675__A1 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15464__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14522__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14095__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13631__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14009__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13924__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13833__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13743__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13632__A1 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15212__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14792__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14370__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13635__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13745__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13636__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15032__I (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14610__I (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14187__I (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13746__I (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13638__I (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13639__A3 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__A3 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A3 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A3 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A3 (.I(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15356__I (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14936__I (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14514__I (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13641__I (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__I (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13929__A1 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13840__A1 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13749__A1 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13643__A1 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A1 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15037__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14615__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14192__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13751__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13646__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13647__A2 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A2 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A2 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A2 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15039__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14617__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14194__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13753__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13649__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13650__A3 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A3 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A3 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A3 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A3 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13653__A1 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13934__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13845__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13756__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13653__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A3 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15376__I (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13655__I (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__I (.I(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14956__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14534__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14107__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13656__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A1 (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14026__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13940__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13849__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13762__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13663__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15364__I (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14944__I (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13757__I (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13658__I (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__I (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13661__I (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13659__A2 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__I (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A1 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13848__A2 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13761__A2 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13662__A2 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15130__I (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14708__I (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14286__I (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13850__I (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13665__I (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13763__A1 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13668__A1 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A2 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A2 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A2 (.I(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15553__I (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14298__I (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13851__I (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13677__I (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13667__I (.I(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13763__B (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13668__B (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15385__I (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13673__I (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__I (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14965__I (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14543__I (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14116__I (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13674__I (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A3 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14031__A3 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13945__A3 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13857__A3 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13767__A3 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13675__A3 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13678__A1 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A2 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13678__A3 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__B (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__B (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__B (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__B (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15387__I (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13679__I (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__I (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14967__I (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14545__I (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14118__I (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13680__I (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__B (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14032__B (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13946__B (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13858__B (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13768__B (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13681__B (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14033__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13947__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13859__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13769__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13683__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13686__A1 (.I(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14052__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13964__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13874__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13783__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13697__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15246__A2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15162__A2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13884__A2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13793__A2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13706__A2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14072__A3 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13986__A3 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13899__A3 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13811__A3 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13718__A3 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13720__A2 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13768__A1 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14076__A1 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13993__A1 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13903__A1 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13815__A1 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13723__A1 (.I(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14080__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13997__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13911__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13819__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13728__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14081__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13998__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13912__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13820__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13730__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14084__A1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14001__A1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13916__A1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13823__A1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13734__A1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14091__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14006__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13921__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13830__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13740__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14099__A3 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14012__A3 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13927__A3 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13838__A3 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13747__A3 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13749__A2 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12023__A1 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14103__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14018__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13931__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13842__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13752__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14104__A3 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14019__A3 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13932__A3 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13843__A3 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13754__A3 (.I(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13756__A1 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13766__A1 (.I(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15043__I (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14621__I (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14198__I (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13758__I (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__I (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14108__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14023__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13935__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13846__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13759__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15394__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15225__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15142__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13863__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13774__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15494__I (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15072__I (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14650__I (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14227__I (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13789__I (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14141__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14058__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13969__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13881__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13790__A1 (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14145__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14062__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13975__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13885__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13795__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15504__I (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15082__I (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14660__I (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14237__I (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13800__I (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14149__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14066__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13980__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13891__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13801__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14152__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14069__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13983__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13896__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13805__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15236__I (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14666__I (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14243__I (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13807__I (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__I (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14154__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14071__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13985__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13898__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13810__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14153__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14070__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13984__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13897__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13809__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13858__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13817__A1 (.I(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13832__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14176__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14086__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14003__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13918__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14175__A1 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14085__A1 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14002__A1 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13917__A1 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13826__A1 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15538__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15116__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14694__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14272__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13836__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14186__A2 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14098__A2 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14011__A2 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13926__A2 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13837__A2 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13844__A2 (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13845__A1 (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14203__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14112__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14027__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13941__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13853__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15131__I (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14709__I (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14287__I (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13951__I (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13852__I (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14203__B (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14112__B (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14027__B (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13941__B (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13853__B (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14214__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14126__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14040__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13953__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13865__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14218__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14130__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14047__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13957__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13870__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14312__I (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13877__I (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A3 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A3 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14224__A3 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14138__A3 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14054__A3 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13966__A3 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13878__A3 (.I(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15586__I (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15164__I (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14744__I (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14322__I (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13887__I (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14234__A1 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14146__A1 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14063__A1 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13976__A1 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13888__A1 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14240__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14151__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14068__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13982__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13895__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14239__A1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14150__A1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14067__A1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13981__A1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13894__A1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13946__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15604__I (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15182__I (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14762__I (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14340__I (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13906__I (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14253__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14164__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14078__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13995__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13907__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15606__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15184__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14764__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14342__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13909__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14254__A2 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14165__A2 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14079__A2 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13996__A2 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13910__A2 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14257__B (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14171__B (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14082__B (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13999__B (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13914__B (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13915__A2 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15358__I (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14938__I (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13938__I (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__I (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__I (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14284__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14201__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14110__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14025__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13939__A2 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13944__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14213__A2 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14125__A2 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14039__A2 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13952__A2 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A3 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13967__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14308__A2 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14220__A2 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14132__A2 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14050__A2 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13960__A2 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14309__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14221__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14133__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14051__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13962__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14311__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14223__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14137__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14053__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13965__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14318__A2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14230__A2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14143__A2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14060__A2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13972__A2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14231__A2 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14144__A2 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14061__A2 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13974__A2 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__A2 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14324__B (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14235__B (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14147__B (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14064__B (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13978__B (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14418__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13989__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__B (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A3 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A3 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14336__A3 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14249__A3 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14159__A3 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14074__A3 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13990__A3 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14032__A1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14337__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14250__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14160__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14075__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13992__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15284__I (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14864__I (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14442__I (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14014__I (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__I (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14362__A1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14276__A1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14190__A1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14101__A1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14016__A1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14018__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14030__A2 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14380__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14295__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14210__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14122__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14035__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14382__A2 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14297__A2 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14212__A2 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14124__A2 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14038__A2 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14385__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14302__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14215__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14127__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14042__A1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15313__I (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14893__I (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14471__I (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14044__I (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__I (.I(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14386__B (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14303__B (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14216__B (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14128__B (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14045__B (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14055__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14390__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14307__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14219__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14131__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14049__A1 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14055__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14399__A1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14315__A1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14226__A1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14140__A1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14057__A1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14083__A1 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14433__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14352__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14265__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14177__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14088__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14434__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14353__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14266__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14180__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14090__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14436__A3 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14355__A3 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14268__A3 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14182__A3 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14093__A3 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14438__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14357__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14270__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14184__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14096__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14115__A1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14454__A1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14372__A1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14285__A1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14202__A1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14111__A1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14115__A2 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14459__A3 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14377__A3 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14292__A3 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14207__A3 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14117__A3 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14460__B (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14378__B (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14293__B (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14208__B (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14119__B (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14461__A1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14379__A1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14294__A1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14209__A1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14121__A1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14125__A1 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15403__I (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14983__I (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14561__I (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14135__I (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__I (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14479__A1 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14395__A1 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14310__A1 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14222__A1 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14136__A1 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14139__A2 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14157__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15424__I (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15003__I (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14581__I (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14156__I (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__I (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14499__A3 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14416__A3 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14334__A3 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14247__A3 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14157__A3 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14158__A2 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14208__A1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14503__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14422__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14338__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14251__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14162__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14172__A1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15434__I (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15013__I (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14591__I (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14167__I (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__I (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14507__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14426__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14344__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14255__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14168__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14508__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14427__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14345__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14256__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14170__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14172__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14511__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14430__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14349__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14259__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14174__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15445__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15024__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14602__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14179__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14518__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14435__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14354__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14267__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14181__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14526__A3 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14441__A3 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14360__A3 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14274__A3 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14188__A3 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14193__A1 (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A1 (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14530__A2 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14446__A2 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14364__A2 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14278__A2 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14193__A2 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14531__A3 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14447__A3 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14365__A3 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14279__A3 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14195__A3 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14206__A1 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14535__A1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14451__A1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14368__A1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14282__A1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14199__A1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14206__A2 (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14212__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14213__A1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14225__A2 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14567__A1 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14485__A1 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14400__A1 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14316__A1 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14228__A1 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14571__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14489__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14405__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14321__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14233__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14575__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14493__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14410__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14326__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14238__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14578__A1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14496__A1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14413__A1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14331__A1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14242__A1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14580__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14498__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14415__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14333__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14246__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14579__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14497__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14414__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14332__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14245__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14248__A2 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14249__A2 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14258__A1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14258__A2 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15527__I (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15105__I (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14683__I (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14261__I (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__I (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14600__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14513__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14432__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14351__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14264__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14599__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14512__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14431__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14350__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14263__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14268__A1 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14609__A2 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14525__A2 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14440__A2 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14359__A2 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14273__A2 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14281__A1 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14291__A1 (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14626__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14539__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14455__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14373__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14288__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14626__B (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14539__B (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14455__B (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14373__B (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14288__B (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14289__A2 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14291__A2 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14636__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14552__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14467__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14383__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14299__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14637__A1 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14553__A1 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14468__A1 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14384__A1 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14301__A1 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14641__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14557__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14474__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14388__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14306__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14647__A3 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14564__A3 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14481__A3 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14397__A3 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14313__A3 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14654__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14570__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14488__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14404__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14320__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14657__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14572__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14490__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14406__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14323__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14663__A2 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14577__A2 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14495__A2 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14412__A2 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14330__A2 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14662__A1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14576__A1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14494__A1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14411__A1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14329__A1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14335__A2 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14378__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14676__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14589__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14505__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14424__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14341__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14677__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14590__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14506__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14425__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14343__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14680__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14595__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14509__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14428__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14347__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14356__A1 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14367__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14376__A1 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14706__A2 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14624__A2 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14537__A2 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14453__A2 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14371__A2 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14376__A2 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14730__A2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14643__A2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14559__A2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14477__A2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14391__A2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14731__A1 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14644__A1 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14560__A1 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14478__A1 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14393__A1 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14733__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14646__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14563__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14480__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14396__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14740__A2 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14653__A2 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14569__A2 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14487__A2 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14403__A2 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14746__B (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14658__B (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14573__B (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14491__B (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14408__B (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14758__A3 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14672__A3 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14584__A3 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14501__A3 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14419__A3 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14460__A1 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14759__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14673__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14585__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14502__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14421__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14784__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14698__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14613__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14528__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14444__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14789__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14703__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14620__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14533__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14450__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14458__A1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14458__A2 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14802__A1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14717__A1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14633__A1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14549__A1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14463__A1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14804__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14719__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14635__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14551__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14466__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14807__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14724__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14638__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14554__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14470__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14808__B (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14725__B (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14639__B (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14555__B (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14472__B (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14812__A1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14729__A1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14642__A1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14558__A1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14476__A1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14821__A1 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14737__A1 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14649__A1 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14566__A1 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14484__A1 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14546__A1 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14855__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14774__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14687__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14601__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14515__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14856__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14775__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14688__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14603__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14517__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14858__A3 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14777__A3 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14690__A3 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14605__A3 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14520__A3 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14860__A1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14779__A1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14692__A1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14607__A1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14523__A1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14542__A1 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14876__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14794__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14707__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14625__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14538__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14881__A3 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14799__A3 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14714__A3 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14630__A3 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14544__A3 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14882__B (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14800__B (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14715__B (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14631__B (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14546__B (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14883__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14801__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14716__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14632__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14548__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14901__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14817__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14732__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14645__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14562__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14582__A1 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14921__A3 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14838__A3 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14756__A3 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14670__A3 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14582__A3 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14631__A1 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14925__A1 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14844__A1 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14760__A1 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14674__A1 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14587__A1 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14929__A1 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14848__A1 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14766__A1 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14678__A1 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14592__A1 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14930__A1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14849__A1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14767__A1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14679__A1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14594__A1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14933__A1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14852__A1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14771__A1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14682__A1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14598__A1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14940__A2 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14857__A2 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14776__A2 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14689__A2 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14604__A2 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14948__A3 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14863__A3 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14782__A3 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14696__A3 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14611__A3 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14952__A2 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14868__A2 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14786__A2 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14700__A2 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14616__A2 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14953__A3 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14869__A3 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14787__A3 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14701__A3 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14618__A3 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14629__A1 (.I(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14957__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14873__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14790__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14704__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14622__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14989__A1 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14907__A1 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14822__A1 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14738__A1 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14651__A1 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14993__A1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14911__A1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14827__A1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14743__A1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14656__A1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14997__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14915__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14832__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14748__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14661__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14670__A1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15000__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14918__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14835__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14753__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14665__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15002__A2 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14920__A2 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14837__A2 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14755__A2 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14669__A2 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15001__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14919__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14836__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14754__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14668__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14715__A1 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15022__A2 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14935__A2 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14854__A2 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14773__A2 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14686__A2 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15021__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14934__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14853__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14772__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14685__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15031__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14947__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14862__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14781__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14695__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14713__A1 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15048__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14961__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14877__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14795__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14710__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15048__B (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14961__B (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14877__B (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14795__B (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14710__B (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15058__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14974__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14889__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14805__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14721__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15059__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14975__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14890__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14806__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14723__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15063__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14979__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14896__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14810__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14728__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15069__A3 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14986__A3 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14903__A3 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14819__A3 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14735__A3 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15076__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14992__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14910__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14826__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14742__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15079__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14994__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14912__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14828__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14745__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15085__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14999__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14917__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14834__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14752__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15084__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14998__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14916__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14833__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14751__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14758__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14800__A1 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15098__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15011__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14927__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14846__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14763__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15099__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15012__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14928__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14847__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14765__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15102__B (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__B (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14931__B (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14850__B (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14769__B (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14784__A2 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12053__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14798__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15128__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15046__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14959__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14875__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14793__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14820__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15151__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15065__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14981__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14899__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14813__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15152__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15066__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14982__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14900__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14815__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15154__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15068__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14985__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14902__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14818__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15161__A2 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15075__A2 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14991__A2 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14909__A2 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14825__A2 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15166__B (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15080__B (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14995__B (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14913__B (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14830__B (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15178__A3 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15094__A3 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15006__A3 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14923__A3 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14841__A3 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14882__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15179__A1 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15095__A1 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15007__A1 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14924__A1 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14843__A1 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15204__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15120__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15035__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14950__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14866__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15209__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15125__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15042__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14955__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14872__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14880__A1 (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15222__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15139__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15055__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14971__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14885__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15224__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15141__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15057__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14973__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14888__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15227__A1 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15145__A1 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15060__A1 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14976__A1 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14892__A1 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15228__B (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15146__B (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15061__B (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14977__B (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14894__B (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15232__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15150__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15064__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14980__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14898__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15241__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15158__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15071__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14988__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14906__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14968__A1 (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15275__A1 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15194__A1 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15109__A1 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15023__A1 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14937__A1 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15276__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15195__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15110__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15025__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14939__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15278__A3 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15197__A3 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15112__A3 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15027__A3 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14942__A3 (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14966__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15280__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15199__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15114__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15029__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14945__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14954__A2 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14964__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15296__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15214__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15129__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15047__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14960__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15301__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15219__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15136__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15052__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14966__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15302__B (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15220__B (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15137__B (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15053__B (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14968__B (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15303__A1 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15221__A1 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15138__A1 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15054__A1 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14970__A1 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15321__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15237__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15153__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15067__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14984__A1 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15341__A3 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15258__A3 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15176__A3 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15092__A3 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15004__A3 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15053__A1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15345__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15264__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15180__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15096__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15009__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15349__A1 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15268__A1 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15186__A1 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15100__A1 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15014__A1 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15350__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15269__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15187__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15101__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15016__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15353__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15272__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15191__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15104__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15020__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15027__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15360__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15277__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15196__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15111__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15026__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15368__A3 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15283__A3 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15202__A3 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15118__A3 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15033__A3 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15372__A2 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15288__A2 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15206__A2 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15122__A2 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15038__A2 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15373__A3 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15289__A3 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15207__A3 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15123__A3 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15040__A3 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15051__A1 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15377__A1 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15293__A1 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15210__A1 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15126__A1 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15044__A1 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15070__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15409__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15327__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15242__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15159__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15073__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15414__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15331__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15247__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15163__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15078__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15418__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15335__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15252__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15168__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15083__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15421__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15338__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15255__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15173__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15087__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15423__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15340__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15257__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15175__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15091__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15422__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15339__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15256__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15174__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15090__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15137__A1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15113__A1 (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15443__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15355__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15274__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15193__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15108__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15442__A1 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15354__A1 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15273__A1 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15192__A1 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15107__A1 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15452__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15367__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15282__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15201__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15117__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15135__A1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15469__A1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15381__A1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15297__A1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15215__A1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15132__A1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15469__B (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15381__B (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15297__B (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15215__B (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15132__B (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15481__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15395__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15310__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15226__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15144__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15485__A1 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15399__A1 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15316__A1 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15230__A1 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15149__A1 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15491__A3 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15406__A3 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15323__A3 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15239__A3 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15156__A3 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15167__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15501__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15415__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15332__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15248__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15165__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15507__A2 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15420__A2 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15337__A2 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15254__A2 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15172__A2 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15506__A1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15419__A1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15336__A1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15253__A1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15171__A1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15177__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15220__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15520__A2 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15432__A2 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15347__A2 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15266__A2 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15183__A2 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15521__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15433__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15348__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15267__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15185__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15524__B (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15438__B (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15351__B (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15270__B (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15189__B (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15198__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15218__A1 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15550__A2 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15467__A2 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15379__A2 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15295__A2 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15213__A2 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15573__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15487__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15401__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15319__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15233__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15574__A1 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15488__A1 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15402__A1 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15320__A1 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15235__A1 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15576__A2 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15490__A2 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15405__A2 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15322__A2 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15238__A2 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15583__A2 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15497__A2 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15411__A2 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15329__A2 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15245__A2 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15588__B (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15502__B (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15416__B (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15333__B (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15250__B (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15259__A2 (.I(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15600__A3 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15516__A3 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15427__A3 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15343__A3 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15261__A3 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15302__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15601__A1 (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15517__A1 (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15428__A1 (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15344__A1 (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15263__A1 (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15279__A1 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15542__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15456__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15370__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15286__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15547__A2 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15463__A2 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15375__A2 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15292__A2 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A2 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15300__A1 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15561__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15476__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15391__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15305__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15563__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15478__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15393__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15308__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15567__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15482__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15396__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15312__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15568__B (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15483__B (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15397__B (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15314__B (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__B (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15572__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15486__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15400__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15318__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15323__A1 (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15580__A1 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15493__A1 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15408__A1 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15326__A1 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A1 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15388__A1 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15531__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15444__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15357__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15532__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15446__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15359__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15534__A3 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15448__A3 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15362__A3 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A3 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A3 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15386__A1 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15536__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15450__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15365__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15384__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15551__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15468__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15380__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15384__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15558__A3 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15473__A3 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15386__A3 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A3 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A3 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15559__B (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15474__B (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15388__B (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__B (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__B (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15560__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15475__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15390__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15575__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15489__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15404__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15498__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15413__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15598__A3 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15514__A3 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15425__A3 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A3 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A3 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15474__A1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15602__A1 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15518__A1 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15430__A1 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A1 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A1 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15608__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15522__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15435__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15609__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15523__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15437__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15526__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15441__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15533__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15447__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15473__A1 (.I(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15540__A3 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15454__A3 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A3 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A3 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A3 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15472__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15548__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15465__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15472__A2 (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15480__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15516__A1 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15581__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15495__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15585__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15500__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15590__A1 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15505__A1 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A1 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A1 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A1 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15595__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15509__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15597__A2 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15513__A2 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A2 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A2 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15596__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15512__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A1 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15514__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15515__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15559__A1 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15530__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15529__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A1 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15558__A1 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15539__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15557__A1 (.I(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15555__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15554__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15554__B (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__B (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__B (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__B (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__B (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15569__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15566__A1 (.I(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__A1 (.I(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A1 (.I(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A1 (.I(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15571__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15573__A1 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15578__A2 (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15578__A3 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A3 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A3 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A3 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A3 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15587__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15594__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15593__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15599__A2 (.I(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15605__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15607__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A2 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15611__B (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__B (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__B (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__B (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__B (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A1 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__A1 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A3 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A2 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A2 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A2 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A2 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__A2 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A1 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A1 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A1 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A1 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A1 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A1 (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A3 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A3 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A3 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A3 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A3 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A1 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A1 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A1 (.I(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__A1 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A2 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A1 (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A1 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__B (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__B (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__B (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__B (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__B (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A1 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A1 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__A1 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A1 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A3 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A3 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A3 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A3 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A3 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A1 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A1 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A1 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A1 (.I(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A3 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A3 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A3 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A3 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__A3 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A2 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__B (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__B (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__B (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__B (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__B (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A2 (.I(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A3 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A3 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__A3 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A3 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A3 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A1 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A1 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A1 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A1 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A2 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A2 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A2 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A3 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A3 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A3 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A3 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A3 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A3 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A3 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A3 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A3 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A3 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A1 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A2 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A3 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__A2 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A2 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A2 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A2 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__A1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A2 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A2 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A1 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A1 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A1 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A1 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A1 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A2 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A2 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A2 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A2 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A1 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A1 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A2 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__I (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__I (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__I (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__I (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__I (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__I (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__I (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__I (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__I (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__I (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__I (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__I (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__I (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__I (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__I (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A1 (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__I (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__I (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__I (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__I (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12287__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__I (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__I (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__B (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__B (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__I (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__I (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__I (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__B (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__B (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__B (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__B (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A1 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A1 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__I (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__I (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__I (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__I (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__I (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__I (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__I (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__I (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__I (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__I (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__A1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__I (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__I (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__I (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__I (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13311__A2 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12176__A2 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__I (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__B (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__B (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__I (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__I (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__B (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__B (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__B (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__B (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__B (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__I (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__I (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__I (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__I (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__I (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__I (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12719__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__I (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__I (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__B (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__B (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__I (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__I (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__I (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__B (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__B (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__B (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__B (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__B (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__I (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__I (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__I (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__I (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__I (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__I (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__I (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__I (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__I (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__I (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__I (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__I (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__I (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__I (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__I (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__I (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__I (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__I (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__I (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__I (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A2 (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13040__A2 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__A2 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__I (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__I (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__B (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__B (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__B (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__B (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__B (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__A1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__I (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__I (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__I (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__I (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__I (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__I (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__I (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__I (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__I (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__I (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__A1 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A1 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A1 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__I (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__I (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__I (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__I (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__I (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__I (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__I (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__I (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__I (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__I (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__A1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__A1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13231__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13151__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__I (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__I (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__B (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__B (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__I (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__I (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__I (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__B (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__B (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__B (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__B (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__B (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A1 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A1 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A1 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A1 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__I (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__I (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__I (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__I (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__I (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__A1 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A1 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A1 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__I (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__I (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__I (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__I (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__I (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13391__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11664__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__I (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__B (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__I (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__I (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__B (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__I (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__I (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__I (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__I (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__I (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__I (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__I (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__I (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__I (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__I (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__I (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__I (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__I (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__I (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__I (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__A1 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A1 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A1 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A1 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A1 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__I (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__I (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__I (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__I (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__I (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11855__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__I (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__I (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__I (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__B (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__B (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__B (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__B (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__B (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A1 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09655__I (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__I (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__I (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__I (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__I (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__I (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__I (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__I (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__I (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__I (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__I (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__I (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12799__A2 (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12095__A2 (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__I (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__I (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__I (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__I (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A2 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__I (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__I (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__I (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__I (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__B (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__B (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__I (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__I (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__I (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__B (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__B (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__B (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__B (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__B (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__B (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__B (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__B (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__B (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__B (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__A2 (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__B (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__I (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__I (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__B (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__I (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__B (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__B (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__B (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__B (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__I (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__I (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__I (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__I (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__I (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A1 (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A1 (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12527__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12447__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__B (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__B (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__B (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__B (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__B (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A1 (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__B (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__B (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__B (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__B (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__B (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__B (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__B (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__I (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__I (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__I (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__B (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__B (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__B (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__B (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__B (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__B (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__B (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__B (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__B (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__B (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A1 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A1 (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A1 (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__B (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__B (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__B (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__B (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__B (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__B (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__B (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__B (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__B (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__B (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A2 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A1 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__B (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__B (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__B (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__B (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__B (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A1 (.I(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A1 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A1 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12367__A1 (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A2 (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__I (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__I (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__I (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__B (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__B (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__B (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__B (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__B (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__A2 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__I (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__I (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__I (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__B (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__B (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__B (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__B (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__B (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A1 (.I(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__B (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__B (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__B (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__B (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__B (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__B (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__B (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__B (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__B (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__B (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A2 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A1 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__B (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__B (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__B (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__B (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__B (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__I (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__I (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__I (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__I (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__I (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__B (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__B (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__B (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__B (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__B (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__B (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__B (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__B (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__B (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__B (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__I (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__I (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__I (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__I (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__I (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A1 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A1 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A1 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A1 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__I (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__I (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__I (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__I (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__I (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A1 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A1 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A1 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A1 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A2 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__B (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__B (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__B (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__B (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__B (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__B (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__B (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__B (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__B (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__B (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A2 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__B (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__B (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__B (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__B (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__B (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A2 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__B (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__B (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__B (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__B (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__B (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A1 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A1 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A1 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A1 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A1 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__A1 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A2 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__B (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__B (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__B (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__B (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__B (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A2 (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A1 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A2 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A2 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A2 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A2 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A2 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__B (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__B (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__B (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__B (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__B (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A1 (.I(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A1 (.I(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__I (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__I (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__I (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__I (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__I (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__A1 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A1 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A1 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A1 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__I (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__I (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__I (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__I (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__I (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A1 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A1 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A1 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A1 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A1 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__B (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__B (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__B (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__B (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__B (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A1 (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A2 (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A1 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__B (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__B (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__B (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__B (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__B (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A1 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A1 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A1 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A1 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A1 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__B (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__B (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__B (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__B (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__B (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A2 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A1 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A1 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A1 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A1 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__I (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__I (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__I (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__I (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__I (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A1 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A1 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A1 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__B (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__B (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__B (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__B (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__B (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A1 (.I(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A2 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A1 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A1 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__A1 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A1 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A1 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A1 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A1 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A1 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A1 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A1 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__B (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__B (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__B (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__B (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__B (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__A1 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A1 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A1 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A1 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A1 (.I(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A1 (.I(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A2 (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A1 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A1 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A1 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A1 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A1 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__B (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__B (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__B (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__B (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__B (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A2 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__A2 (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A1 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A1 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A1 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A1 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A1 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A1 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A1 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A1 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A1 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__A2 (.I(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A1 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A1 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A1 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A1 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A1 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A1 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A1 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A1 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A1 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A1 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A1 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A2 (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__A1 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A1 (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A2 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__I (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__I (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__I (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__I (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__B (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__B (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__B (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__B (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__B (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__A1 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__B (.I(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__B (.I(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__B (.I(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__B (.I(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__B (.I(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A1 (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A1 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A1 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A1 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A1 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__B (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__B (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__B (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__B (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__B (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A2 (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A1 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A1 (.I(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A1 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A1 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A1 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A1 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A1 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A1 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A1 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A1 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A1 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A1 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__A1 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A1 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A1 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A1 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A1 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A2 (.I(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A1 (.I(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A1 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A1 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A1 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A1 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A1 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A1 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A2 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A1 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A1 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A1 (.I(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A2 (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__A1 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__A1 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A1 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A1 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A1 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A1 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A1 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A1 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A1 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A1 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A1 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A1 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A1 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A1 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A2 (.I(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A2 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__B (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__B (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__B (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__B (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__B (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__A2 (.I(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__A1 (.I(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A1 (.I(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A1 (.I(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A1 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A1 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__B (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__B (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__B (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__B (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__B (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A1 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A1 (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A1 (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A1 (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A1 (.I(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A1 (.I(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A1 (.I(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A1 (.I(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A1 (.I(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A1 (.I(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A1 (.I(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A1 (.I(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A2 (.I(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A1 (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A1 (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A1 (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A1 (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A1 (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A2 (.I(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__B (.I(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__B (.I(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__B (.I(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__B (.I(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__B (.I(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__A1 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A1 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A1 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A1 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A1 (.I(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A1 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A1 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A2 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A1 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A1 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A1 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A1 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__A1 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__B (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__B (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__B (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__B (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__B (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__B (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__B (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__B (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__B (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__B (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A2 (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A2 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A1 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A1 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A1 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A2 (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A1 (.I(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A1 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A1 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A2 (.I(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A2 (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A1 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__A1 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A1 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__A1 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__A1 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A1 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A1 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A1 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A1 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A1 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A1 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A1 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A1 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A1 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A1 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__A1 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A1 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A1 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A2 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A1 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A1 (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A2 (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A1 (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A1 (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__A1 (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__A1 (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A1 (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A1 (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A1 (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A2 (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A2 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A1 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A1 (.I(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A1 (.I(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A1 (.I(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A1 (.I(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A1 (.I(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__A1 (.I(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A1 (.I(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A1 (.I(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A1 (.I(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__A1 (.I(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__A1 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A1 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A1 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__A1 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A1 (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A1 (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A1 (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A1 (.I(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__B (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__B (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__B (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__B (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__B (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A2 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A2 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A1 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A1 (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A1 (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A1 (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__A1 (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A2 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A2 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A2 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A2 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A2 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__B (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__B (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__B (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__B (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__B (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A1 (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A1 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A2 (.I(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__A1 (.I(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A1 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A1 (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A1 (.I(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A1 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A1 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__A1 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A1 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A1 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A1 (.I(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A2 (.I(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A1 (.I(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A1 (.I(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A1 (.I(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A1 (.I(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A1 (.I(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A1 (.I(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A1 (.I(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__B (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__B (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__B (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__B (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__B (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A1 (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__A1 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A1 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A1 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A1 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A1 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A1 (.I(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A1 (.I(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A1 (.I(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A1 (.I(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__A1 (.I(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A1 (.I(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A1 (.I(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__A1 (.I(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A2 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A1 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A1 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A1 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A1 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A1 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A1 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A1 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A1 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A1 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A1 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A1 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A1 (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A1 (.I(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__A1 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A1 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__A1 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A1 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A1 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A1 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A1 (.I(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__A1 (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A1 (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A1 (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A1 (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A2 (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A2 (.I(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__A1 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A1 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A1 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A1 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A1 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A2 (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A1 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A2 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A1 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A1 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A1 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A1 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A1 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A2 (.I(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A1 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__A1 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A1 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A1 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A2 (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A1 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A1 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A1 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A1 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A1 (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A1 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A1 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__A1 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A1 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A2 (.I(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A1 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A2 (.I(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A1 (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A1 (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A1 (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A1 (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A1 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__A1 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__A1 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A1 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A1 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A2 (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__A2 (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A2 (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A2 (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A2 (.I(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A1 (.I(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A1 (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A1 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A1 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A1 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A1 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A1 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__A1 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A1 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A1 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A1 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A1 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A1 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A2 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A2 (.I(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A1 (.I(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A1 (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A1 (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A1 (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__A1 (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A1 (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A1 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A1 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__A1 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__A1 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A1 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A2 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__A1 (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__A2 (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__A1 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A1 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__A1 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A1 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A1 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A1 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A1 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A1 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__A1 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A1 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A2 (.I(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A1 (.I(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A1 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A1 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A1 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A1 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A1 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A1 (.I(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A1 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__A1 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A1 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A1 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A1 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A2 (.I(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__A1 (.I(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A2 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A2 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A1 (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A1 (.I(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__A2 (.I(_05884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__A1 (.I(_05885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A2 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__A1 (.I(_05906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A1 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__A2 (.I(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A1 (.I(_05930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A1 (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A1 (.I(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A2 (.I(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__A2 (.I(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A1 (.I(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A1 (.I(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A1 (.I(_05996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A2 (.I(_06003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__I (.I(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12175__I (.I(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11663__I (.I(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__I (.I(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__I (.I(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A1 (.I(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A1 (.I(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A1 (.I(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A1 (.I(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11855__A1 (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__A1 (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A1 (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__A1 (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__I (.I(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__I (.I(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__I (.I(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__I (.I(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A1 (.I(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A1 (.I(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A1 (.I(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__A1 (.I(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__I (.I(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__I (.I(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__I (.I(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__I (.I(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__I (.I(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__I (.I(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A2 (.I(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A2 (.I(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A1 (.I(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A1 (.I(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A1 (.I(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12615__I (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12183__I (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__I (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__I (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__I (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A1 (.I(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A1 (.I(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A1 (.I(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A1 (.I(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A1 (.I(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12618__I (.I(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12186__I (.I(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__I (.I(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__I (.I(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__I (.I(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A1 (.I(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__A1 (.I(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A1 (.I(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A1 (.I(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12621__I (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12189__I (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__I (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__I (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__I (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A1 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__A1 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A1 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A1 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A1 (.I(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A1 (.I(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A1 (.I(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A1 (.I(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A1 (.I(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13057__I (.I(_06044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__I (.I(_06044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12625__I (.I(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12193__I (.I(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11681__I (.I(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__I (.I(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__I (.I(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__A1 (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A1 (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A1 (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A1 (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__A1 (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13060__I (.I(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__I (.I(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12628__I (.I(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12196__I (.I(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__I (.I(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__I (.I(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__I (.I(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A1 (.I(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A1 (.I(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__I (.I(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__I (.I(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__I (.I(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__I (.I(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__I (.I(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A2 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A2 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A2 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A2 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13065__I (.I(_06054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__I (.I(_06054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12633__I (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__I (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11689__I (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__I (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__I (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A1 (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__A1 (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A1 (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A1 (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A1 (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13068__I (.I(_06058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__I (.I(_06058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12636__I (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12204__I (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11692__I (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__I (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__I (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__A1 (.I(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__A1 (.I(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A1 (.I(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A1 (.I(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13071__I (.I(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__I (.I(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12639__I (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12207__I (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__I (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__I (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__I (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A1 (.I(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A1 (.I(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A1 (.I(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A1 (.I(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A1 (.I(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13075__I (.I(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__I (.I(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12643__I (.I(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12211__I (.I(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__I (.I(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__I (.I(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__I (.I(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A1 (.I(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A1 (.I(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A1 (.I(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A1 (.I(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A1 (.I(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12646__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12214__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11702__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A1 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A1 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A1 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A1 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A1 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A2 (.I(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A2 (.I(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A2 (.I(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__A2 (.I(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A2 (.I(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12650__I (.I(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12218__I (.I(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11706__I (.I(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__I (.I(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__I (.I(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A1 (.I(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A1 (.I(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__A1 (.I(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__A1 (.I(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12653__I (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12221__I (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__I (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__I (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__I (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__A1 (.I(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A1 (.I(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A1 (.I(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A1 (.I(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A1 (.I(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12656__I (.I(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__I (.I(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__I (.I(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__I (.I(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__I (.I(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A1 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__A1 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A1 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A1 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A1 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A1 (.I(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A1 (.I(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__A1 (.I(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A1 (.I(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12660__I (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12228__I (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11716__I (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__I (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__I (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A1 (.I(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__A1 (.I(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A1 (.I(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A1 (.I(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A1 (.I(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12663__I (.I(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12231__I (.I(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__I (.I(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__I (.I(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__I (.I(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A1 (.I(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A1 (.I(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A1 (.I(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A1 (.I(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A2 (.I(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A2 (.I(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A2 (.I(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A2 (.I(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A2 (.I(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12667__I (.I(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12235__I (.I(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11723__I (.I(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__I (.I(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__I (.I(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A1 (.I(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A1 (.I(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A1 (.I(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A1 (.I(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12670__I (.I(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__I (.I(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11726__I (.I(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I (.I(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__I (.I(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A1 (.I(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A1 (.I(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A1 (.I(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A1 (.I(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12673__I (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12241__I (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11729__I (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11297__I (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__I (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__A1 (.I(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A1 (.I(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A1 (.I(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A1 (.I(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A1 (.I(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A1 (.I(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A1 (.I(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A1 (.I(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A1 (.I(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A1 (.I(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12677__I (.I(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12245__I (.I(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11733__I (.I(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__I (.I(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__I (.I(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A1 (.I(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A1 (.I(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A1 (.I(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A1 (.I(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13112__I (.I(_06115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__I (.I(_06115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12680__I (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12248__I (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11736__I (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__I (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__I (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A1 (.I(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__A1 (.I(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__A1 (.I(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A1 (.I(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A1 (.I(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__A2 (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__A2 (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A2 (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A2 (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A2 (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13116__I (.I(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__I (.I(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12684__I (.I(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12252__I (.I(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11740__I (.I(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__I (.I(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__I (.I(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__A1 (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A1 (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A1 (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A1 (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A1 (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13119__I (.I(_06124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__I (.I(_06124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__I (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12255__I (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11743__I (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__I (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__I (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A1 (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A1 (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A1 (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A1 (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A1 (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__I (.I(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12258__I (.I(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11746__I (.I(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__I (.I(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__I (.I(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__A1 (.I(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A1 (.I(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A1 (.I(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__A1 (.I(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A1 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A1 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__A1 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A1 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__A1 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12694__I (.I(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12262__I (.I(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__I (.I(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__I (.I(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__I (.I(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A1 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A1 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A1 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A1 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__A1 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13129__I (.I(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__I (.I(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12697__I (.I(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12265__I (.I(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11753__I (.I(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__I (.I(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__I (.I(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__A1 (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A1 (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A1 (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A1 (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12701__I (.I(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12269__I (.I(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11757__I (.I(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__I (.I(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__I (.I(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A1 (.I(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__A1 (.I(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A1 (.I(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A1 (.I(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A1 (.I(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13136__I (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__I (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12704__I (.I(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12272__I (.I(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11760__I (.I(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__I (.I(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__I (.I(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__A1 (.I(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__A1 (.I(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__A1 (.I(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A1 (.I(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A1 (.I(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__I (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12275__I (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11763__I (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__I (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__I (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A1 (.I(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A1 (.I(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A1 (.I(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A1 (.I(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A1 (.I(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12710__I (.I(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12278__I (.I(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11766__I (.I(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__I (.I(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__I (.I(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__A1 (.I(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__A1 (.I(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A1 (.I(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A1 (.I(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A1 (.I(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12713__I (.I(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12281__I (.I(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11769__I (.I(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__I (.I(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__I (.I(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__A1 (.I(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A1 (.I(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A1 (.I(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A1 (.I(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12716__I (.I(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12284__I (.I(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__I (.I(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__I (.I(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__I (.I(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A1 (.I(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A1 (.I(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A1 (.I(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A1 (.I(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A1 (.I(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__I (.I(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__I (.I(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__I (.I(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__I (.I(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A1 (.I(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A1 (.I(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A1 (.I(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A1 (.I(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__I (.I(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A2 (.I(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A2 (.I(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A2 (.I(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A2 (.I(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A2 (.I(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__I (.I(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__I (.I(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__I (.I(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__I (.I(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__I (.I(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A2 (.I(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A2 (.I(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A1 (.I(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A1 (.I(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A1 (.I(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A1 (.I(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A1 (.I(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A1 (.I(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__A1 (.I(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__I (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__I (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__I (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__I (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__I (.I(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A2 (.I(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A2 (.I(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A2 (.I(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A2 (.I(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A2 (.I(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A1 (.I(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A1 (.I(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A1 (.I(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A1 (.I(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A2 (.I(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A2 (.I(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A2 (.I(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A2 (.I(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A2 (.I(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A1 (.I(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A1 (.I(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A1 (.I(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A1 (.I(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A1 (.I(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A2 (.I(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A2 (.I(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A2 (.I(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A2 (.I(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A2 (.I(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A1 (.I(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A1 (.I(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A1 (.I(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A1 (.I(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A1 (.I(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A2 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A2 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A2 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A2 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A2 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A1 (.I(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A1 (.I(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A1 (.I(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A1 (.I(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A2 (.I(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A2 (.I(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A2 (.I(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A2 (.I(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A2 (.I(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12015__A2 (.I(_06214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__I (.I(_06214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13040__A1 (.I(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12719__A1 (.I(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11664__A1 (.I(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__A1 (.I(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__A2 (.I(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__I (.I(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__I (.I(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__I (.I(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__I (.I(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A1 (.I(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__A1 (.I(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A1 (.I(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A1 (.I(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__I (.I(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A2 (.I(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A2 (.I(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A2 (.I(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A2 (.I(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A2 (.I(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__I (.I(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__I (.I(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__I (.I(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__I (.I(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__I (.I(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A2 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A2 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A1 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__A1 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A1 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A1 (.I(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A1 (.I(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__A1 (.I(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A1 (.I(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A1 (.I(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__I (.I(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__I (.I(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__I (.I(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__I (.I(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__I (.I(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A2 (.I(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A2 (.I(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A2 (.I(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A2 (.I(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A2 (.I(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A1 (.I(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A2 (.I(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A2 (.I(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A2 (.I(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__A2 (.I(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A2 (.I(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__A1 (.I(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__A1 (.I(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A1 (.I(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A1 (.I(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A2 (.I(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A2 (.I(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A2 (.I(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A2 (.I(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A2 (.I(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A1 (.I(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A1 (.I(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A1 (.I(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__A1 (.I(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A2 (.I(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A2 (.I(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A2 (.I(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A2 (.I(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__A2 (.I(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A1 (.I(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A1 (.I(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A1 (.I(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A1 (.I(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__A1 (.I(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A2 (.I(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A2 (.I(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__A2 (.I(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A2 (.I(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A2 (.I(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12095__A1 (.I(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__A1 (.I(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__A1 (.I(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A1 (.I(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A1 (.I(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__I (.I(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__I (.I(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__I (.I(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__I (.I(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__A1 (.I(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A1 (.I(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A1 (.I(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__I (.I(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A2 (.I(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__A2 (.I(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__A2 (.I(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A2 (.I(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A2 (.I(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__I (.I(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__I (.I(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__I (.I(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__I (.I(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__I (.I(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A2 (.I(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A2 (.I(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__A1 (.I(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__A1 (.I(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__A1 (.I(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A1 (.I(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__A1 (.I(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A1 (.I(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A1 (.I(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__I (.I(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__I (.I(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__I (.I(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__I (.I(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__I (.I(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A2 (.I(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A2 (.I(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__A2 (.I(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__A2 (.I(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A2 (.I(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__A1 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A1 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A1 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__A1 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__B (.I(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__A2 (.I(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__A2 (.I(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A2 (.I(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A2 (.I(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A2 (.I(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A1 (.I(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A1 (.I(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__A1 (.I(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A1 (.I(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A1 (.I(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A2 (.I(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A2 (.I(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A2 (.I(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A2 (.I(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A2 (.I(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A1 (.I(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__A1 (.I(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A1 (.I(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A1 (.I(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__A1 (.I(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A2 (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A2 (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A2 (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A2 (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__A2 (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A1 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A1 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__A1 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A1 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A1 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__A2 (.I(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A2 (.I(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__A2 (.I(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__A2 (.I(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A2 (.I(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13391__A1 (.I(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13311__A1 (.I(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__A1 (.I(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__I (.I(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12799__A1 (.I(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__A1 (.I(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12287__A1 (.I(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11935__A1 (.I(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__A1 (.I(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__I (.I(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__I (.I(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__I (.I(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__I (.I(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__A1 (.I(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11227__A1 (.I(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A1 (.I(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__A1 (.I(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__I (.I(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__A2 (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A2 (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A2 (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A2 (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A2 (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__I (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__I (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__I (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__I (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__I (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A2 (.I(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__A2 (.I(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__A1 (.I(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A1 (.I(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__A1 (.I(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A1 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A1 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A1 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__A1 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__I (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__I (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__I (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__I (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__I (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A2 (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A2 (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__A2 (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A2 (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A2 (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A1 (.I(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A1 (.I(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A1 (.I(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A1 (.I(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A1 (.I(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__B (.I(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__B (.I(_06336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A2 (.I(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A2 (.I(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__A2 (.I(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A2 (.I(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A2 (.I(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A1 (.I(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A1 (.I(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A1 (.I(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A1 (.I(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A1 (.I(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A2 (.I(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__A2 (.I(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A2 (.I(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A2 (.I(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A2 (.I(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A1 (.I(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11207__A1 (.I(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A1 (.I(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A1 (.I(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A2 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__A2 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A2 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__A2 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A2 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A1 (.I(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A1 (.I(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A1 (.I(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__A1 (.I(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A1 (.I(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__A2 (.I(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A2 (.I(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__A2 (.I(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A2 (.I(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__A2 (.I(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__A1 (.I(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__A1 (.I(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__A1 (.I(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A1 (.I(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__A1 (.I(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__I (.I(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__I (.I(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__I (.I(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__I (.I(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A1 (.I(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A1 (.I(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A1 (.I(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A1 (.I(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__I (.I(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A2 (.I(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A2 (.I(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A2 (.I(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A2 (.I(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__A2 (.I(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__I (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__I (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__I (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__I (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__I (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A2 (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A2 (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A1 (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A1 (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A1 (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__A1 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__A1 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A1 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A1 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A1 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A1 (.I(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__A1 (.I(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11433__A1 (.I(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A1 (.I(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__A1 (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A1 (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__A1 (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A1 (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A1 (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A1 (.I(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A1 (.I(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A1 (.I(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A1 (.I(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__A1 (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A1 (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__A1 (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A1 (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A1 (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A1 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A1 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A1 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A1 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A1 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__I (.I(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__I (.I(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__I (.I(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__I (.I(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__I (.I(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A2 (.I(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A2 (.I(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A2 (.I(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A2 (.I(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A2 (.I(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A1 (.I(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A1 (.I(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__A1 (.I(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__A1 (.I(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A1 (.I(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__A1 (.I(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__A1 (.I(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__A1 (.I(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A1 (.I(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__A1 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__A1 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__A1 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A1 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A1 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__A1 (.I(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A1 (.I(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A1 (.I(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A1 (.I(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A1 (.I(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__A1 (.I(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__A1 (.I(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A1 (.I(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__A1 (.I(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A1 (.I(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__A1 (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11534__A1 (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__A1 (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A1 (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A1 (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A2 (.I(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__A2 (.I(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A2 (.I(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A2 (.I(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A2 (.I(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A1 (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A1 (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A1 (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__A1 (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__A1 (.I(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A1 (.I(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A1 (.I(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__A1 (.I(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A1 (.I(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__A1 (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A1 (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A1 (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A1 (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__A1 (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__A1 (.I(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__A1 (.I(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A1 (.I(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A1 (.I(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A1 (.I(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A1 (.I(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__A1 (.I(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__A1 (.I(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A1 (.I(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A1 (.I(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A2 (.I(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A2 (.I(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A2 (.I(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A2 (.I(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A2 (.I(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__A1 (.I(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__A1 (.I(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A1 (.I(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A1 (.I(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A1 (.I(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A1 (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11550__A1 (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__A1 (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11390__A1 (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A1 (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__A1 (.I(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__A1 (.I(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__A1 (.I(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A1 (.I(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A1 (.I(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A1 (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A1 (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A1 (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A1 (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A1 (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__A1 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A1 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__A1 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A1 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A1 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__A1 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__A1 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__A1 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A1 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A1 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__A1 (.I(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__A1 (.I(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__A1 (.I(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A1 (.I(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A1 (.I(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A1 (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__A1 (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A1 (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A1 (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__A1 (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__A1 (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A1 (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__A1 (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A1 (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__A1 (.I(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A1 (.I(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__A1 (.I(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__A1 (.I(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A1 (.I(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11647__A1 (.I(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__A1 (.I(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__A1 (.I(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A1 (.I(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11650__A1 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__A1 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__A1 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A1 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A1 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__A2 (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A2 (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__A2 (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A2 (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A2 (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11652__A1 (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A1 (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A1 (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A1 (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A1 (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__A1 (.I(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__A1 (.I(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__A1 (.I(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A1 (.I(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__A1 (.I(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__A1 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__A1 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__A1 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A1 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__A1 (.I(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A1 (.I(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A1 (.I(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A1 (.I(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__A1 (.I(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__A1 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A1 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11500__A1 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A1 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__A1 (.I(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A1 (.I(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__A1 (.I(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A1 (.I(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A1 (.I(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__I (.I(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__I (.I(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__I (.I(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__I (.I(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A1 (.I(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A1 (.I(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A1 (.I(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A1 (.I(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__I (.I(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A2 (.I(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A2 (.I(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A2 (.I(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A2 (.I(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A2 (.I(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__I (.I(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__I (.I(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__I (.I(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__I (.I(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__I (.I(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A2 (.I(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A2 (.I(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A1 (.I(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A1 (.I(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A1 (.I(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__A1 (.I(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__A1 (.I(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A1 (.I(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__A1 (.I(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__A1 (.I(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__I (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__I (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__I (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__I (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__I (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__A2 (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A2 (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__A2 (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__A2 (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A2 (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11377__A1 (.I(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A1 (.I(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A1 (.I(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A1 (.I(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__A1 (.I(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A2 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A2 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__A2 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__A2 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A2 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__A1 (.I(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A1 (.I(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A1 (.I(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A1 (.I(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A1 (.I(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A2 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A2 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11390__A2 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A2 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A2 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A1 (.I(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A1 (.I(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__A1 (.I(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__A1 (.I(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__A1 (.I(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A2 (.I(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__A2 (.I(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A2 (.I(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A2 (.I(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A2 (.I(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A1 (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A1 (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A1 (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__A1 (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A1 (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A2 (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A2 (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A2 (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A2 (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A2 (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11483__I (.I(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__I (.I(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__I (.I(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__I (.I(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__A1 (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__A1 (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__A1 (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A1 (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__I (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__A2 (.I(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__A2 (.I(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11433__A2 (.I(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A2 (.I(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__A2 (.I(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__I (.I(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__I (.I(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11439__I (.I(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__I (.I(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__I (.I(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__A2 (.I(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11500__A2 (.I(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A1 (.I(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__A1 (.I(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__A1 (.I(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__A1 (.I(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__A1 (.I(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__A1 (.I(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A1 (.I(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A1 (.I(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__I (.I(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__I (.I(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__I (.I(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__I (.I(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__I (.I(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A2 (.I(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__A2 (.I(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__A2 (.I(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__A2 (.I(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A2 (.I(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A1 (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A1 (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A1 (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__A1 (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A1 (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A2 (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A2 (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A2 (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A2 (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__A2 (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A1 (.I(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A1 (.I(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__A1 (.I(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__A1 (.I(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__A1 (.I(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__A2 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__A2 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__A2 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A2 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__A2 (.I(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__A1 (.I(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A1 (.I(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__A1 (.I(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__A1 (.I(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__A1 (.I(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__A2 (.I(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A2 (.I(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A2 (.I(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__A2 (.I(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__A2 (.I(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A1 (.I(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11491__A1 (.I(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11489__A1 (.I(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__A1 (.I(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__A1 (.I(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A2 (.I(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__A2 (.I(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__A2 (.I(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A2 (.I(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__A2 (.I(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__I (.I(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__I (.I(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__I (.I(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__I (.I(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11581__A1 (.I(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A1 (.I(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__A1 (.I(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__A1 (.I(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__I (.I(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A2 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A2 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__A2 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__A2 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__A2 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11539__I (.I(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11527__I (.I(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__I (.I(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__I (.I(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__I (.I(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A2 (.I(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A2 (.I(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A1 (.I(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__A1 (.I(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__A1 (.I(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__A1 (.I(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A1 (.I(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__A1 (.I(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__A1 (.I(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__A1 (.I(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__I (.I(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__I (.I(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__I (.I(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__I (.I(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__I (.I(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__A2 (.I(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__A2 (.I(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__A2 (.I(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A2 (.I(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A2 (.I(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__A1 (.I(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A1 (.I(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__A1 (.I(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__A1 (.I(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__A1 (.I(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__A2 (.I(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A2 (.I(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A2 (.I(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A2 (.I(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11534__A2 (.I(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__A1 (.I(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__A1 (.I(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__A1 (.I(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__A1 (.I(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11540__A1 (.I(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A2 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__A2 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11550__A2 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__A2 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__A2 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A1 (.I(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A1 (.I(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__A1 (.I(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__A1 (.I(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A1 (.I(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__A2 (.I(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__A2 (.I(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__A2 (.I(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__A2 (.I(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__A2 (.I(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__A1 (.I(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A1 (.I(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__A1 (.I(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__A1 (.I(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__A1 (.I(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A2 (.I(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__A2 (.I(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__A2 (.I(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A2 (.I(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__A2 (.I(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__I (.I(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11631__I (.I(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11586__I (.I(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__I (.I(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11661__A1 (.I(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__A1 (.I(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11657__A1 (.I(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__A1 (.I(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__I (.I(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__A2 (.I(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__A2 (.I(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A2 (.I(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__A2 (.I(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__A2 (.I(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__I (.I(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__I (.I(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11599__I (.I(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__I (.I(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__I (.I(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__A2 (.I(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__A2 (.I(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__A1 (.I(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11590__A1 (.I(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__A1 (.I(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11603__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11597__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11648__I (.I(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11636__I (.I(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__I (.I(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__I (.I(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__I (.I(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__A2 (.I(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__A2 (.I(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A2 (.I(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A2 (.I(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A2 (.I(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__A1 (.I(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__A1 (.I(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__A1 (.I(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__A1 (.I(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__A1 (.I(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__A2 (.I(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__A2 (.I(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__A2 (.I(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A2 (.I(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__A2 (.I(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11629__A1 (.I(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__A1 (.I(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11625__A1 (.I(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__A1 (.I(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__A1 (.I(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__A2 (.I(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__A2 (.I(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A2 (.I(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__A2 (.I(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A2 (.I(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11641__A1 (.I(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11639__A1 (.I(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11637__A1 (.I(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__A1 (.I(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__A1 (.I(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11647__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11649__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__A2 (.I(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__A2 (.I(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__A2 (.I(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11652__A2 (.I(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11650__A2 (.I(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12101__A1 (.I(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__A1 (.I(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11861__A1 (.I(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11781__A1 (.I(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A1 (.I(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11747__I (.I(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11730__I (.I(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__I (.I(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__I (.I(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__A1 (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__A1 (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11767__A1 (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__A1 (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__I (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__A2 (.I(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__A2 (.I(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__A2 (.I(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__A2 (.I(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A2 (.I(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__I (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__I (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__I (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__I (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__I (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11774__A2 (.I(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11771__A2 (.I(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__A1 (.I(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__A1 (.I(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__A1 (.I(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12103__A1 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11943__A1 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__A1 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__A1 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__A1 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12105__A1 (.I(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__A1 (.I(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__A1 (.I(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11785__A1 (.I(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__A1 (.I(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12108__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11948__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11868__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__A1 (.I(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11690__A1 (.I(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__A1 (.I(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__A1 (.I(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__A1 (.I(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12110__A1 (.I(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__A1 (.I(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11870__A1 (.I(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11790__A1 (.I(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__A1 (.I(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12114__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11954__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11874__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11754__I (.I(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11737__I (.I(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__I (.I(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__I (.I(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11686__I (.I(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__A2 (.I(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__A2 (.I(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11694__A2 (.I(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11691__A2 (.I(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__A2 (.I(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12116__A1 (.I(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11956__A1 (.I(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__A1 (.I(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__A1 (.I(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11691__A1 (.I(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12118__A1 (.I(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11958__A1 (.I(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__A1 (.I(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__A1 (.I(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11694__A1 (.I(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12121__A1 (.I(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11961__A1 (.I(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11881__A1 (.I(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11801__A1 (.I(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__A1 (.I(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11710__A1 (.I(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__A1 (.I(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11704__A1 (.I(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__A1 (.I(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__A1 (.I(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__A1 (.I(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__A1 (.I(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11883__A1 (.I(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__A1 (.I(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__A1 (.I(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12126__A1 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11966__A1 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11886__A1 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11806__A1 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__A1 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11708__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12128__A1 (.I(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11968__A1 (.I(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11888__A1 (.I(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__A1 (.I(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11708__A1 (.I(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12130__A1 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11970__A1 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11890__A1 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11810__A1 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__A1 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12133__A1 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__A1 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11893__A1 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__A1 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A1 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__A1 (.I(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11724__A1 (.I(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__A1 (.I(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__A1 (.I(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A1 (.I(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12135__A1 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__A1 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11895__A1 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__A1 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__A1 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12138__A1 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__A1 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11898__A1 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__A1 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11722__A1 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__A2 (.I(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11732__A2 (.I(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11728__A2 (.I(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11725__A2 (.I(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11722__A2 (.I(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12140__A1 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__A1 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11900__A1 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11820__A1 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11725__A1 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12142__A1 (.I(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__A1 (.I(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__A1 (.I(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11822__A1 (.I(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11728__A1 (.I(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12145__A1 (.I(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11985__A1 (.I(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__A1 (.I(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11825__A1 (.I(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11732__A1 (.I(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11744__A1 (.I(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__A1 (.I(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11738__A1 (.I(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11734__A1 (.I(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__A1 (.I(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12147__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11987__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12150__A1 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__A1 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11910__A1 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11830__A1 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__A1 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__A2 (.I(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11749__A2 (.I(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__A2 (.I(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__A2 (.I(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__A2 (.I(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12152__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11832__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12154__A1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11994__A1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11914__A1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__A1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__A1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12157__A1 (.I(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11997__A1 (.I(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__A1 (.I(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__A1 (.I(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11749__A1 (.I(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__A1 (.I(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__A1 (.I(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11755__A1 (.I(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11751__A1 (.I(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__A1 (.I(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12159__A1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__A1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__A1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__A1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12162__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11922__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11768__A2 (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11765__A2 (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11762__A2 (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11759__A2 (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__A2 (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12164__A1 (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__A1 (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__A1 (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11844__A1 (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11759__A1 (.I(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12166__A1 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12006__A1 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__A1 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11846__A1 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11762__A1 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12168__A1 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12008__A1 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__A1 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__A1 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11765__A1 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12170__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12010__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11850__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11768__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12172__A1 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12012__A1 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__A1 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11852__A1 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11771__A1 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12174__A1 (.I(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12014__A1 (.I(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__A1 (.I(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__A1 (.I(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11774__A1 (.I(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__I (.I(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11823__I (.I(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11778__I (.I(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11776__I (.I(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11853__A1 (.I(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11851__A1 (.I(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11849__A1 (.I(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11847__A1 (.I(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11777__I (.I(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11790__A2 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__A2 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11785__A2 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__A2 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11781__A2 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11811__I (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11799__I (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__I (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11786__I (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11779__I (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__A2 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11852__A2 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__A1 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__A1 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11780__A1 (.I(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11797__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11795__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11789__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11840__I (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11828__I (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__I (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__I (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11792__I (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11801__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11809__A1 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__A1 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__A1 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11802__A1 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__A1 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__A2 (.I(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__A2 (.I(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11810__A2 (.I(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__A2 (.I(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11806__A2 (.I(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11821__A1 (.I(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__A1 (.I(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__A1 (.I(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__A1 (.I(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11812__A1 (.I(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11825__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11822__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11820__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__A1 (.I(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__A1 (.I(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11829__A1 (.I(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11826__A1 (.I(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11824__A1 (.I(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A2 (.I(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__A2 (.I(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__A2 (.I(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11832__A2 (.I(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11830__A2 (.I(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__A1 (.I(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11843__A1 (.I(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11841__A1 (.I(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__A1 (.I(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11836__A1 (.I(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11850__A2 (.I(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__A2 (.I(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11846__A2 (.I(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11844__A2 (.I(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__A2 (.I(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11915__I (.I(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11903__I (.I(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11858__I (.I(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11856__I (.I(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__A1 (.I(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__A1 (.I(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__A1 (.I(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11927__A1 (.I(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__I (.I(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11870__A2 (.I(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11868__A2 (.I(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__A2 (.I(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__A2 (.I(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11861__A2 (.I(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11891__I (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11879__I (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__I (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11866__I (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11859__I (.I(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__A2 (.I(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__A2 (.I(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11864__A1 (.I(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__A1 (.I(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11860__A1 (.I(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11920__I (.I(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11908__I (.I(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11896__I (.I(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11884__I (.I(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11872__I (.I(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11883__A2 (.I(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11881__A2 (.I(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__A2 (.I(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__A2 (.I(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11874__A2 (.I(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11889__A1 (.I(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11887__A1 (.I(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11885__A1 (.I(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11882__A1 (.I(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11880__A1 (.I(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11895__A2 (.I(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11893__A2 (.I(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11890__A2 (.I(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11888__A2 (.I(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11886__A2 (.I(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__A1 (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11899__A1 (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11897__A1 (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11894__A1 (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11892__A1 (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__A2 (.I(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__A2 (.I(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__A2 (.I(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11900__A2 (.I(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11898__A2 (.I(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__A1 (.I(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11911__A1 (.I(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__A1 (.I(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11906__A1 (.I(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11904__A1 (.I(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__A2 (.I(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__A2 (.I(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11914__A2 (.I(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__A2 (.I(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11910__A2 (.I(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11925__A1 (.I(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11923__A1 (.I(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11921__A1 (.I(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11918__A1 (.I(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11916__A1 (.I(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__A2 (.I(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__A2 (.I(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__A2 (.I(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__A2 (.I(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11922__A2 (.I(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11995__I (.I(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11983__I (.I(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11938__I (.I(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11936__I (.I(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12013__A1 (.I(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12011__A1 (.I(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__A1 (.I(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__A1 (.I(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__I (.I(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__A2 (.I(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11948__A2 (.I(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__A2 (.I(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11943__A2 (.I(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__A2 (.I(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11971__I (.I(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11959__I (.I(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11951__I (.I(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__I (.I(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11939__I (.I(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12014__A2 (.I(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12012__A2 (.I(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11944__A1 (.I(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11942__A1 (.I(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__A1 (.I(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__A1 (.I(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__A1 (.I(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__A1 (.I(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11949__A1 (.I(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11947__A1 (.I(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12000__I (.I(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11988__I (.I(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11976__I (.I(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__I (.I(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11952__I (.I(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11954__B (.I(_06827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__A1 (.I(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11967__A1 (.I(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11965__A1 (.I(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__A1 (.I(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__A1 (.I(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__B (.I(_06832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__A2 (.I(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__A2 (.I(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11970__A2 (.I(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11968__A2 (.I(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11966__A2 (.I(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11981__A1 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11979__A1 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__A1 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11974__A1 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11972__A1 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11987__A2 (.I(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11985__A2 (.I(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__A2 (.I(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__A2 (.I(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__A2 (.I(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__A1 (.I(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11991__A1 (.I(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__A1 (.I(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11986__A1 (.I(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11984__A1 (.I(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__A2 (.I(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11997__A2 (.I(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11994__A2 (.I(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__A2 (.I(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__A2 (.I(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12005__A1 (.I(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12003__A1 (.I(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__A1 (.I(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__A1 (.I(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11996__A1 (.I(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12010__A2 (.I(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12008__A2 (.I(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12006__A2 (.I(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__A2 (.I(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__A2 (.I(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12075__I (.I(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12063__I (.I(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__I (.I(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12016__I (.I(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12093__A1 (.I(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12091__A1 (.I(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12089__A1 (.I(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12087__A1 (.I(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12017__I (.I(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12030__A2 (.I(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12028__A2 (.I(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12025__A2 (.I(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12023__A2 (.I(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12021__A2 (.I(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12051__I (.I(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__I (.I(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__I (.I(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12026__I (.I(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12019__I (.I(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12094__A2 (.I(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12092__A2 (.I(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12024__A1 (.I(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12022__A1 (.I(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__A1 (.I(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__A1 (.I(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__A1 (.I(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12033__A1 (.I(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__A1 (.I(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__A1 (.I(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12080__I (.I(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12068__I (.I(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12056__I (.I(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12044__I (.I(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__I (.I(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12043__A2 (.I(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__A2 (.I(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12038__A2 (.I(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12036__A2 (.I(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12034__A2 (.I(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12034__B (.I(_06875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12049__A1 (.I(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__A1 (.I(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A1 (.I(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12042__A1 (.I(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__A1 (.I(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12055__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12053__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12050__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12048__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12046__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12061__A1 (.I(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12059__A1 (.I(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12057__A1 (.I(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12054__A1 (.I(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12052__A1 (.I(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12067__A2 (.I(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12065__A2 (.I(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12062__A2 (.I(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12060__A2 (.I(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12058__A2 (.I(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12073__A1 (.I(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12071__A1 (.I(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12069__A1 (.I(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12066__A1 (.I(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12064__A1 (.I(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12065__B (.I(_06893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__A2 (.I(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12077__A2 (.I(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12074__A2 (.I(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12072__A2 (.I(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12070__A2 (.I(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12090__A2 (.I(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12088__A2 (.I(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12086__A2 (.I(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12084__A2 (.I(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12082__A2 (.I(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12082__B (.I(_06903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12084__B (.I(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12086__B (.I(_06905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12155__I (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12143__I (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12098__I (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12096__I (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12173__A1 (.I(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12171__A1 (.I(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12169__A1 (.I(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12167__A1 (.I(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12097__I (.I(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12110__A2 (.I(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12108__A2 (.I(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12105__A2 (.I(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12103__A2 (.I(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12101__A2 (.I(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12131__I (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12119__I (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12111__I (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12106__I (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12099__I (.I(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12174__A2 (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12172__A2 (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__A1 (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12102__A1 (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12100__A1 (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__A1 (.I(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12115__A1 (.I(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12113__A1 (.I(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12109__A1 (.I(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__A1 (.I(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12160__I (.I(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12148__I (.I(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12136__I (.I(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12124__I (.I(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12112__I (.I(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__A2 (.I(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12121__A2 (.I(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12118__A2 (.I(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12116__A2 (.I(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12114__A2 (.I(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12129__A1 (.I(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12127__A1 (.I(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12125__A1 (.I(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12122__A1 (.I(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12120__A1 (.I(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12135__A2 (.I(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12133__A2 (.I(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12130__A2 (.I(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12128__A2 (.I(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12126__A2 (.I(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12141__A1 (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12139__A1 (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12137__A1 (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12134__A1 (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12132__A1 (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12147__A2 (.I(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12145__A2 (.I(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12142__A2 (.I(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12140__A2 (.I(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12138__A2 (.I(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__A1 (.I(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12151__A1 (.I(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__A1 (.I(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12146__A1 (.I(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12144__A1 (.I(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12159__A2 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12157__A2 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12154__A2 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12152__A2 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12150__A2 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12165__A1 (.I(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12163__A1 (.I(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12161__A1 (.I(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12158__A1 (.I(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12156__A1 (.I(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12170__A2 (.I(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12168__A2 (.I(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12166__A2 (.I(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12164__A2 (.I(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12162__A2 (.I(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12533__A1 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12453__A1 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12373__A1 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12293__A1 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12182__A1 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12259__I (.I(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__I (.I(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12179__I (.I(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12177__I (.I(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12285__A1 (.I(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12282__A1 (.I(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12279__A1 (.I(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12276__A1 (.I(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12178__I (.I(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__A2 (.I(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12192__A2 (.I(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__A2 (.I(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__A2 (.I(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12182__A2 (.I(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12225__I (.I(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12208__I (.I(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12197__I (.I(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12190__I (.I(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__I (.I(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12286__A2 (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12283__A2 (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12187__A1 (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__A1 (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12181__A1 (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12535__A1 (.I(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12455__A1 (.I(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12375__A1 (.I(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12295__A1 (.I(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__A1 (.I(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12537__A1 (.I(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12457__A1 (.I(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12377__A1 (.I(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12297__A1 (.I(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__A1 (.I(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12540__A1 (.I(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__A1 (.I(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12380__A1 (.I(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12300__A1 (.I(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12192__A1 (.I(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12205__A1 (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12202__A1 (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12199__A1 (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12194__A1 (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12191__A1 (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12542__A1 (.I(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12462__A1 (.I(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12382__A1 (.I(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12302__A1 (.I(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__A1 (.I(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12546__A1 (.I(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12466__A1 (.I(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12386__A1 (.I(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12306__A1 (.I(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__A1 (.I(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12266__I (.I(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12249__I (.I(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12232__I (.I(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__I (.I(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12198__I (.I(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__A2 (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12210__A2 (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__A2 (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12203__A2 (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__A2 (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12548__A1 (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12468__A1 (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12388__A1 (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12308__A1 (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12203__A1 (.I(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12550__A1 (.I(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12470__A1 (.I(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12390__A1 (.I(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12310__A1 (.I(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__A1 (.I(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12553__A1 (.I(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12473__A1 (.I(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12393__A1 (.I(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12313__A1 (.I(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12210__A1 (.I(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12222__A1 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12219__A1 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12216__A1 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12212__A1 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A1 (.I(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12555__A1 (.I(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__A1 (.I(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12395__A1 (.I(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12315__A1 (.I(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__A1 (.I(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__A1 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12478__A1 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12398__A1 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__A1 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12217__A1 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__A2 (.I(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12227__A2 (.I(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__A2 (.I(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12220__A2 (.I(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12217__A2 (.I(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12560__A1 (.I(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12480__A1 (.I(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12400__A1 (.I(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12320__A1 (.I(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12220__A1 (.I(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12562__A1 (.I(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__A1 (.I(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12402__A1 (.I(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12322__A1 (.I(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__A1 (.I(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12565__A1 (.I(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12485__A1 (.I(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12405__A1 (.I(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12325__A1 (.I(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12227__A1 (.I(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__A1 (.I(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12236__A1 (.I(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__A1 (.I(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__A1 (.I(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12226__A1 (.I(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12567__A1 (.I(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12487__A1 (.I(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12407__A1 (.I(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12327__A1 (.I(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__A1 (.I(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12570__A1 (.I(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12490__A1 (.I(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12410__A1 (.I(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12330__A1 (.I(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12234__A1 (.I(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12247__A2 (.I(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12244__A2 (.I(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12240__A2 (.I(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__A2 (.I(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12234__A2 (.I(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12572__A1 (.I(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12492__A1 (.I(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12412__A1 (.I(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12332__A1 (.I(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__A1 (.I(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12574__A1 (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12494__A1 (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12414__A1 (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12334__A1 (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12240__A1 (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12577__A1 (.I(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12497__A1 (.I(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12417__A1 (.I(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12337__A1 (.I(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12244__A1 (.I(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12256__A1 (.I(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12253__A1 (.I(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12250__A1 (.I(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12246__A1 (.I(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12243__A1 (.I(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12579__A1 (.I(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12499__A1 (.I(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12419__A1 (.I(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12339__A1 (.I(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12247__A1 (.I(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__A1 (.I(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12502__A1 (.I(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12422__A1 (.I(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12342__A1 (.I(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12251__A1 (.I(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12264__A2 (.I(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12261__A2 (.I(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12257__A2 (.I(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12254__A2 (.I(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12251__A2 (.I(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12584__A1 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12504__A1 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12424__A1 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12344__A1 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12254__A1 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12586__A1 (.I(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12506__A1 (.I(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12426__A1 (.I(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12346__A1 (.I(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12257__A1 (.I(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12589__A1 (.I(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12509__A1 (.I(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12429__A1 (.I(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12349__A1 (.I(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12261__A1 (.I(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12273__A1 (.I(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12270__A1 (.I(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12267__A1 (.I(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12263__A1 (.I(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12260__A1 (.I(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12591__A1 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12511__A1 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12431__A1 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12351__A1 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12264__A1 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12594__A1 (.I(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12514__A1 (.I(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12434__A1 (.I(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12354__A1 (.I(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12268__A1 (.I(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12280__A2 (.I(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12277__A2 (.I(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12274__A2 (.I(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12271__A2 (.I(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12268__A2 (.I(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12516__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12436__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12356__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12271__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12598__A1 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__A1 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12438__A1 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12358__A1 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12274__A1 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12600__A1 (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A1 (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12440__A1 (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12360__A1 (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12277__A1 (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__A1 (.I(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12522__A1 (.I(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12442__A1 (.I(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12362__A1 (.I(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12280__A1 (.I(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12604__A1 (.I(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12524__A1 (.I(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12444__A1 (.I(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12364__A1 (.I(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12283__A1 (.I(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12606__A1 (.I(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__A1 (.I(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12446__A1 (.I(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12366__A1 (.I(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12286__A1 (.I(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12347__I (.I(_07038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12335__I (.I(_07038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12290__I (.I(_07038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12288__I (.I(_07038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__A1 (.I(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12363__A1 (.I(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12361__A1 (.I(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12359__A1 (.I(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12289__I (.I(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12302__A2 (.I(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12300__A2 (.I(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12297__A2 (.I(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12295__A2 (.I(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12293__A2 (.I(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12323__I (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12311__I (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12303__I (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12298__I (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12291__I (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12366__A2 (.I(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12364__A2 (.I(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12296__A1 (.I(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12294__A1 (.I(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__A1 (.I(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__A1 (.I(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12307__A1 (.I(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12305__A1 (.I(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12301__A1 (.I(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12299__A1 (.I(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12352__I (.I(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12340__I (.I(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12328__I (.I(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12316__I (.I(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12304__I (.I(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12315__A2 (.I(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12313__A2 (.I(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12310__A2 (.I(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12308__A2 (.I(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12306__A2 (.I(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12321__A1 (.I(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12319__A1 (.I(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12317__A1 (.I(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12314__A1 (.I(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12312__A1 (.I(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12327__A2 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12325__A2 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12322__A2 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12320__A2 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__A2 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12333__A1 (.I(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12331__A1 (.I(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12329__A1 (.I(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12326__A1 (.I(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12324__A1 (.I(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12339__A2 (.I(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12337__A2 (.I(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12334__A2 (.I(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12332__A2 (.I(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12330__A2 (.I(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12345__A1 (.I(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12343__A1 (.I(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12341__A1 (.I(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12338__A1 (.I(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12336__A1 (.I(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12351__A2 (.I(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12349__A2 (.I(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12346__A2 (.I(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12344__A2 (.I(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12342__A2 (.I(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12357__A1 (.I(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12355__A1 (.I(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12353__A1 (.I(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12350__A1 (.I(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12348__A1 (.I(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12362__A2 (.I(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12360__A2 (.I(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12358__A2 (.I(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12356__A2 (.I(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12354__A2 (.I(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12427__I (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12415__I (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__I (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12368__I (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12445__A1 (.I(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__A1 (.I(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12441__A1 (.I(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12439__A1 (.I(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12369__I (.I(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12382__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12380__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12377__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12375__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12373__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12403__I (.I(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12391__I (.I(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12383__I (.I(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12378__I (.I(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12371__I (.I(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12446__A2 (.I(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12444__A2 (.I(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12376__A1 (.I(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12374__A1 (.I(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12372__A1 (.I(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12389__A1 (.I(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12387__A1 (.I(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12385__A1 (.I(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12381__A1 (.I(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12379__A1 (.I(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12432__I (.I(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12420__I (.I(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12408__I (.I(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12396__I (.I(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12384__I (.I(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12395__A2 (.I(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12393__A2 (.I(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12390__A2 (.I(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12388__A2 (.I(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12386__A2 (.I(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12401__A1 (.I(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12399__A1 (.I(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12397__A1 (.I(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12394__A1 (.I(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12392__A1 (.I(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12407__A2 (.I(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12405__A2 (.I(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12402__A2 (.I(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12400__A2 (.I(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12398__A2 (.I(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12413__A1 (.I(_07109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12411__A1 (.I(_07109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12409__A1 (.I(_07109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12406__A1 (.I(_07109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12404__A1 (.I(_07109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12419__A2 (.I(_07112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12417__A2 (.I(_07112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12414__A2 (.I(_07112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12412__A2 (.I(_07112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12410__A2 (.I(_07112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12425__A1 (.I(_07116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12423__A1 (.I(_07116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12421__A1 (.I(_07116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12418__A1 (.I(_07116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12416__A1 (.I(_07116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12431__A2 (.I(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12429__A2 (.I(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12426__A2 (.I(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12424__A2 (.I(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12422__A2 (.I(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12437__A1 (.I(_07123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12435__A1 (.I(_07123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12433__A1 (.I(_07123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12430__A1 (.I(_07123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12428__A1 (.I(_07123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12442__A2 (.I(_07126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12440__A2 (.I(_07126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12438__A2 (.I(_07126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12436__A2 (.I(_07126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12434__A2 (.I(_07126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12507__I (.I(_07134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12495__I (.I(_07134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12450__I (.I(_07134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12448__I (.I(_07134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__A1 (.I(_07135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12523__A1 (.I(_07135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12521__A1 (.I(_07135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12519__A1 (.I(_07135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12449__I (.I(_07135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12462__A2 (.I(_07136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__A2 (.I(_07136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12457__A2 (.I(_07136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12455__A2 (.I(_07136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12453__A2 (.I(_07136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12483__I (.I(_07137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12471__I (.I(_07137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12463__I (.I(_07137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12458__I (.I(_07137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12451__I (.I(_07137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__A2 (.I(_07138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12524__A2 (.I(_07138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12456__A1 (.I(_07138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12454__A1 (.I(_07138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12452__A1 (.I(_07138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12469__A1 (.I(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12467__A1 (.I(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12465__A1 (.I(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__A1 (.I(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12459__A1 (.I(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12512__I (.I(_07145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12500__I (.I(_07145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12488__I (.I(_07145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12476__I (.I(_07145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12464__I (.I(_07145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__A2 (.I(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12473__A2 (.I(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12470__A2 (.I(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12468__A2 (.I(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12466__A2 (.I(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__A1 (.I(_07150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12479__A1 (.I(_07150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12477__A1 (.I(_07150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12474__A1 (.I(_07150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12472__A1 (.I(_07150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12487__A2 (.I(_07153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12485__A2 (.I(_07153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__A2 (.I(_07153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12480__A2 (.I(_07153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12478__A2 (.I(_07153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12493__A1 (.I(_07157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12491__A1 (.I(_07157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__A1 (.I(_07157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12486__A1 (.I(_07157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12484__A1 (.I(_07157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12499__A2 (.I(_07160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12497__A2 (.I(_07160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12494__A2 (.I(_07160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12492__A2 (.I(_07160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12490__A2 (.I(_07160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12505__A1 (.I(_07164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12503__A1 (.I(_07164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12501__A1 (.I(_07164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12498__A1 (.I(_07164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12496__A1 (.I(_07164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12511__A2 (.I(_07167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12509__A2 (.I(_07167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12506__A2 (.I(_07167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12504__A2 (.I(_07167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12502__A2 (.I(_07167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__A1 (.I(_07171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12515__A1 (.I(_07171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12513__A1 (.I(_07171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12510__A1 (.I(_07171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12508__A1 (.I(_07171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12522__A2 (.I(_07174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A2 (.I(_07174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__A2 (.I(_07174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12516__A2 (.I(_07174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12514__A2 (.I(_07174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12587__I (.I(_07182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12575__I (.I(_07182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12530__I (.I(_07182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12528__I (.I(_07182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12605__A1 (.I(_07183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__A1 (.I(_07183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12601__A1 (.I(_07183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12599__A1 (.I(_07183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12529__I (.I(_07183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12542__A2 (.I(_07184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12540__A2 (.I(_07184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12537__A2 (.I(_07184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12535__A2 (.I(_07184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12533__A2 (.I(_07184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12563__I (.I(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12551__I (.I(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12543__I (.I(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12538__I (.I(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12531__I (.I(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12606__A2 (.I(_07186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12604__A2 (.I(_07186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__A1 (.I(_07186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__A1 (.I(_07186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12532__A1 (.I(_07186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12549__A1 (.I(_07190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__A1 (.I(_07190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12545__A1 (.I(_07190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12541__A1 (.I(_07190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12539__A1 (.I(_07190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12592__I (.I(_07193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12580__I (.I(_07193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12568__I (.I(_07193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12556__I (.I(_07193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12544__I (.I(_07193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12555__A2 (.I(_07194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12553__A2 (.I(_07194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12550__A2 (.I(_07194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12548__A2 (.I(_07194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12546__A2 (.I(_07194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12561__A1 (.I(_07198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12559__A1 (.I(_07198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12557__A1 (.I(_07198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12554__A1 (.I(_07198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12552__A1 (.I(_07198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12567__A2 (.I(_07201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12565__A2 (.I(_07201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12562__A2 (.I(_07201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12560__A2 (.I(_07201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__A2 (.I(_07201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12573__A1 (.I(_07205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12571__A1 (.I(_07205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12569__A1 (.I(_07205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12566__A1 (.I(_07205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12564__A1 (.I(_07205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12579__A2 (.I(_07208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12577__A2 (.I(_07208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12574__A2 (.I(_07208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12572__A2 (.I(_07208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12570__A2 (.I(_07208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12585__A1 (.I(_07212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__A1 (.I(_07212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12581__A1 (.I(_07212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12578__A1 (.I(_07212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12576__A1 (.I(_07212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12591__A2 (.I(_07215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12589__A2 (.I(_07215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12586__A2 (.I(_07215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12584__A2 (.I(_07215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__A2 (.I(_07215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12597__A1 (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12595__A1 (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12593__A1 (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12590__A1 (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12588__A1 (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__A2 (.I(_07222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12600__A2 (.I(_07222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12598__A2 (.I(_07222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__A2 (.I(_07222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12594__A2 (.I(_07222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12965__A1 (.I(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12885__A1 (.I(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12805__A1 (.I(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12725__A1 (.I(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12614__A1 (.I(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__I (.I(_07231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12674__I (.I(_07231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12611__I (.I(_07231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12609__I (.I(_07231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12717__A1 (.I(_07232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12714__A1 (.I(_07232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12711__A1 (.I(_07232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12708__A1 (.I(_07232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12610__I (.I(_07232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12627__A2 (.I(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12624__A2 (.I(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12620__A2 (.I(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12617__A2 (.I(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12614__A2 (.I(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12657__I (.I(_07234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12640__I (.I(_07234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12629__I (.I(_07234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12622__I (.I(_07234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__I (.I(_07234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12718__A2 (.I(_07235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12715__A2 (.I(_07235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12619__A1 (.I(_07235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12616__A1 (.I(_07235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12613__A1 (.I(_07235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12967__A1 (.I(_07237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12887__A1 (.I(_07237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12807__A1 (.I(_07237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12727__A1 (.I(_07237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12617__A1 (.I(_07237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12969__A1 (.I(_07239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12889__A1 (.I(_07239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12809__A1 (.I(_07239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__A1 (.I(_07239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12620__A1 (.I(_07239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12972__A1 (.I(_07241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12892__A1 (.I(_07241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12812__A1 (.I(_07241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12732__A1 (.I(_07241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12624__A1 (.I(_07241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__A1 (.I(_07242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12634__A1 (.I(_07242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12631__A1 (.I(_07242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__A1 (.I(_07242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__A1 (.I(_07242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12974__A1 (.I(_07244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12894__A1 (.I(_07244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12814__A1 (.I(_07244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12734__A1 (.I(_07244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12627__A1 (.I(_07244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12978__A1 (.I(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12898__A1 (.I(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12818__A1 (.I(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12738__A1 (.I(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12632__A1 (.I(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12698__I (.I(_07247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12681__I (.I(_07247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12664__I (.I(_07247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12647__I (.I(_07247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12630__I (.I(_07247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12645__A2 (.I(_07248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__A2 (.I(_07248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12638__A2 (.I(_07248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12635__A2 (.I(_07248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12632__A2 (.I(_07248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12980__A1 (.I(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12900__A1 (.I(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12820__A1 (.I(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12740__A1 (.I(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12635__A1 (.I(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12982__A1 (.I(_07252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12902__A1 (.I(_07252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__A1 (.I(_07252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12742__A1 (.I(_07252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12638__A1 (.I(_07252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12985__A1 (.I(_07254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12905__A1 (.I(_07254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12825__A1 (.I(_07254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12745__A1 (.I(_07254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__A1 (.I(_07254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12654__A1 (.I(_07255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12651__A1 (.I(_07255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12648__A1 (.I(_07255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12644__A1 (.I(_07255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12641__A1 (.I(_07255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12987__A1 (.I(_07257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12907__A1 (.I(_07257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12827__A1 (.I(_07257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12747__A1 (.I(_07257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12645__A1 (.I(_07257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12990__A1 (.I(_07259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__A1 (.I(_07259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12830__A1 (.I(_07259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12750__A1 (.I(_07259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12649__A1 (.I(_07259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12662__A2 (.I(_07260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12659__A2 (.I(_07260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12655__A2 (.I(_07260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12652__A2 (.I(_07260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12649__A2 (.I(_07260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12992__A1 (.I(_07262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12912__A1 (.I(_07262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12832__A1 (.I(_07262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12752__A1 (.I(_07262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12652__A1 (.I(_07262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12994__A1 (.I(_07264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12914__A1 (.I(_07264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12834__A1 (.I(_07264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12754__A1 (.I(_07264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12655__A1 (.I(_07264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12997__A1 (.I(_07266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12917__A1 (.I(_07266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12837__A1 (.I(_07266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12757__A1 (.I(_07266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12659__A1 (.I(_07266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12671__A1 (.I(_07267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12668__A1 (.I(_07267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12665__A1 (.I(_07267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__A1 (.I(_07267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12658__A1 (.I(_07267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12999__A1 (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12919__A1 (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12839__A1 (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12759__A1 (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12662__A1 (.I(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13002__A1 (.I(_07271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12922__A1 (.I(_07271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12842__A1 (.I(_07271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12762__A1 (.I(_07271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12666__A1 (.I(_07271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12679__A2 (.I(_07272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12676__A2 (.I(_07272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12672__A2 (.I(_07272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12669__A2 (.I(_07272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12666__A2 (.I(_07272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13004__A1 (.I(_07274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12924__A1 (.I(_07274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12844__A1 (.I(_07274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12764__A1 (.I(_07274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12669__A1 (.I(_07274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13006__A1 (.I(_07276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12926__A1 (.I(_07276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12846__A1 (.I(_07276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12766__A1 (.I(_07276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12672__A1 (.I(_07276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13009__A1 (.I(_07278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12929__A1 (.I(_07278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12849__A1 (.I(_07278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12769__A1 (.I(_07278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12676__A1 (.I(_07278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12688__A1 (.I(_07279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12685__A1 (.I(_07279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12682__A1 (.I(_07279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12678__A1 (.I(_07279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12675__A1 (.I(_07279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13011__A1 (.I(_07281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12931__A1 (.I(_07281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12851__A1 (.I(_07281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12771__A1 (.I(_07281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12679__A1 (.I(_07281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13014__A1 (.I(_07283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12934__A1 (.I(_07283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12854__A1 (.I(_07283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12774__A1 (.I(_07283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12683__A1 (.I(_07283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12696__A2 (.I(_07284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12693__A2 (.I(_07284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12689__A2 (.I(_07284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__A2 (.I(_07284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12683__A2 (.I(_07284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13016__A1 (.I(_07286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12936__A1 (.I(_07286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12856__A1 (.I(_07286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12776__A1 (.I(_07286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__A1 (.I(_07286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13018__A1 (.I(_07288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12938__A1 (.I(_07288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12858__A1 (.I(_07288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12778__A1 (.I(_07288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12689__A1 (.I(_07288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13021__A1 (.I(_07290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12941__A1 (.I(_07290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12861__A1 (.I(_07290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12781__A1 (.I(_07290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12693__A1 (.I(_07290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__A1 (.I(_07291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12702__A1 (.I(_07291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12699__A1 (.I(_07291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12695__A1 (.I(_07291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12692__A1 (.I(_07291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13023__A1 (.I(_07293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12943__A1 (.I(_07293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12863__A1 (.I(_07293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12783__A1 (.I(_07293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12696__A1 (.I(_07293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13026__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12946__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12866__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12700__A1 (.I(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12712__A2 (.I(_07296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12709__A2 (.I(_07296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12706__A2 (.I(_07296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__A2 (.I(_07296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12700__A2 (.I(_07296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13028__A1 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12948__A1 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12868__A1 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__A1 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__A1 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13030__A1 (.I(_07300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12950__A1 (.I(_07300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12870__A1 (.I(_07300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12790__A1 (.I(_07300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12706__A1 (.I(_07300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13032__A1 (.I(_07302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12952__A1 (.I(_07302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12872__A1 (.I(_07302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12792__A1 (.I(_07302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12709__A1 (.I(_07302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13034__A1 (.I(_07304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12954__A1 (.I(_07304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12874__A1 (.I(_07304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12794__A1 (.I(_07304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12712__A1 (.I(_07304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13036__A1 (.I(_07306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12956__A1 (.I(_07306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12876__A1 (.I(_07306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12796__A1 (.I(_07306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12715__A1 (.I(_07306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13038__A1 (.I(_07308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12958__A1 (.I(_07308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12878__A1 (.I(_07308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12798__A1 (.I(_07308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12718__A1 (.I(_07308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12779__I (.I(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12767__I (.I(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12722__I (.I(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12720__I (.I(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12797__A1 (.I(_07311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12795__A1 (.I(_07311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12793__A1 (.I(_07311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12791__A1 (.I(_07311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12721__I (.I(_07311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12734__A2 (.I(_07312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12732__A2 (.I(_07312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__A2 (.I(_07312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12727__A2 (.I(_07312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12725__A2 (.I(_07312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12755__I (.I(_07313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12743__I (.I(_07313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12735__I (.I(_07313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12730__I (.I(_07313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12723__I (.I(_07313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12798__A2 (.I(_07314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12796__A2 (.I(_07314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12728__A1 (.I(_07314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12726__A1 (.I(_07314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12724__A1 (.I(_07314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12741__A1 (.I(_07318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12739__A1 (.I(_07318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12737__A1 (.I(_07318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12733__A1 (.I(_07318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12731__A1 (.I(_07318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12784__I (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12772__I (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12760__I (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12748__I (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12736__I (.I(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12747__A2 (.I(_07322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12745__A2 (.I(_07322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12742__A2 (.I(_07322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12740__A2 (.I(_07322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12738__A2 (.I(_07322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12738__B (.I(_07323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12740__B (.I(_07324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12753__A1 (.I(_07326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12751__A1 (.I(_07326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__A1 (.I(_07326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12746__A1 (.I(_07326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12744__A1 (.I(_07326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12759__A2 (.I(_07329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12757__A2 (.I(_07329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12754__A2 (.I(_07329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12752__A2 (.I(_07329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12750__A2 (.I(_07329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12765__A1 (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12763__A1 (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12761__A1 (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12758__A1 (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12756__A1 (.I(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12771__A2 (.I(_07336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12769__A2 (.I(_07336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12766__A2 (.I(_07336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12764__A2 (.I(_07336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12762__A2 (.I(_07336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12777__A1 (.I(_07340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12775__A1 (.I(_07340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12773__A1 (.I(_07340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12770__A1 (.I(_07340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12768__A1 (.I(_07340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12783__A2 (.I(_07343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12781__A2 (.I(_07343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12778__A2 (.I(_07343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12776__A2 (.I(_07343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12774__A2 (.I(_07343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12789__A1 (.I(_07347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12787__A1 (.I(_07347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12785__A1 (.I(_07347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12782__A1 (.I(_07347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12780__A1 (.I(_07347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12794__A2 (.I(_07350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12792__A2 (.I(_07350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12790__A2 (.I(_07350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__A2 (.I(_07350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__A2 (.I(_07350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12859__I (.I(_07358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12847__I (.I(_07358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12802__I (.I(_07358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12800__I (.I(_07358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12877__A1 (.I(_07359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12875__A1 (.I(_07359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12873__A1 (.I(_07359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12871__A1 (.I(_07359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12801__I (.I(_07359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12814__A2 (.I(_07360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12812__A2 (.I(_07360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12809__A2 (.I(_07360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12807__A2 (.I(_07360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12805__A2 (.I(_07360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12835__I (.I(_07361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12823__I (.I(_07361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12815__I (.I(_07361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12810__I (.I(_07361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12803__I (.I(_07361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12878__A2 (.I(_07362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12876__A2 (.I(_07362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12808__A1 (.I(_07362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12806__A1 (.I(_07362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12804__A1 (.I(_07362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12821__A1 (.I(_07366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12819__A1 (.I(_07366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12817__A1 (.I(_07366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12813__A1 (.I(_07366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12811__A1 (.I(_07366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12864__I (.I(_07369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12852__I (.I(_07369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12840__I (.I(_07369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12828__I (.I(_07369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__I (.I(_07369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12827__A2 (.I(_07370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12825__A2 (.I(_07370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__A2 (.I(_07370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12820__A2 (.I(_07370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12818__A2 (.I(_07370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12820__B (.I(_07372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12833__A1 (.I(_07374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12831__A1 (.I(_07374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12829__A1 (.I(_07374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12826__A1 (.I(_07374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12824__A1 (.I(_07374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12839__A2 (.I(_07377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12837__A2 (.I(_07377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12834__A2 (.I(_07377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12832__A2 (.I(_07377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12830__A2 (.I(_07377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__A1 (.I(_07381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12843__A1 (.I(_07381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12841__A1 (.I(_07381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12838__A1 (.I(_07381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12836__A1 (.I(_07381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12851__A2 (.I(_07384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12849__A2 (.I(_07384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12846__A2 (.I(_07384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12844__A2 (.I(_07384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12842__A2 (.I(_07384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12857__A1 (.I(_07388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12855__A1 (.I(_07388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12853__A1 (.I(_07388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12850__A1 (.I(_07388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12848__A1 (.I(_07388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12863__A2 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12861__A2 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12858__A2 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12856__A2 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12854__A2 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__A1 (.I(_07395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12867__A1 (.I(_07395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12865__A1 (.I(_07395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12862__A1 (.I(_07395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12860__A1 (.I(_07395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12874__A2 (.I(_07398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12872__A2 (.I(_07398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12870__A2 (.I(_07398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12868__A2 (.I(_07398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12866__A2 (.I(_07398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12939__I (.I(_07406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12927__I (.I(_07406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12882__I (.I(_07406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12880__I (.I(_07406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12957__A1 (.I(_07407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12955__A1 (.I(_07407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12953__A1 (.I(_07407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12951__A1 (.I(_07407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__I (.I(_07407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12894__A2 (.I(_07408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12892__A2 (.I(_07408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12889__A2 (.I(_07408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12887__A2 (.I(_07408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12885__A2 (.I(_07408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12915__I (.I(_07409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12903__I (.I(_07409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12895__I (.I(_07409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12890__I (.I(_07409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12883__I (.I(_07409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12958__A2 (.I(_07410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12956__A2 (.I(_07410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12888__A1 (.I(_07410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12886__A1 (.I(_07410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12884__A1 (.I(_07410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12901__A1 (.I(_07414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12899__A1 (.I(_07414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12897__A1 (.I(_07414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12893__A1 (.I(_07414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12891__A1 (.I(_07414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12944__I (.I(_07417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12932__I (.I(_07417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12920__I (.I(_07417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__I (.I(_07417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12896__I (.I(_07417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12907__A2 (.I(_07418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12905__A2 (.I(_07418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12902__A2 (.I(_07418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12900__A2 (.I(_07418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12898__A2 (.I(_07418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12898__B (.I(_07419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12913__A1 (.I(_07422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12911__A1 (.I(_07422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__A1 (.I(_07422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12906__A1 (.I(_07422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12904__A1 (.I(_07422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12919__A2 (.I(_07425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12917__A2 (.I(_07425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12914__A2 (.I(_07425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12912__A2 (.I(_07425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__A2 (.I(_07425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12925__A1 (.I(_07429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12923__A1 (.I(_07429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12921__A1 (.I(_07429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12918__A1 (.I(_07429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__A1 (.I(_07429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12931__A2 (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12929__A2 (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12926__A2 (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12924__A2 (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12922__A2 (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12937__A1 (.I(_07436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12935__A1 (.I(_07436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12933__A1 (.I(_07436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12930__A1 (.I(_07436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12928__A1 (.I(_07436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12943__A2 (.I(_07439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12941__A2 (.I(_07439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12938__A2 (.I(_07439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12936__A2 (.I(_07439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12934__A2 (.I(_07439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12949__A1 (.I(_07443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__A1 (.I(_07443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12945__A1 (.I(_07443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12942__A1 (.I(_07443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12940__A1 (.I(_07443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12954__A2 (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12952__A2 (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12950__A2 (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12948__A2 (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12946__A2 (.I(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13019__I (.I(_07454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13007__I (.I(_07454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12962__I (.I(_07454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12960__I (.I(_07454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13037__A1 (.I(_07455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13035__A1 (.I(_07455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13033__A1 (.I(_07455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13031__A1 (.I(_07455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12961__I (.I(_07455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12974__A2 (.I(_07456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12972__A2 (.I(_07456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12969__A2 (.I(_07456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12967__A2 (.I(_07456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12965__A2 (.I(_07456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12995__I (.I(_07457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12983__I (.I(_07457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12975__I (.I(_07457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12970__I (.I(_07457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12963__I (.I(_07457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13038__A2 (.I(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13036__A2 (.I(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12968__A1 (.I(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12966__A1 (.I(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12964__A1 (.I(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12981__A1 (.I(_07462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12979__A1 (.I(_07462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12977__A1 (.I(_07462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12973__A1 (.I(_07462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12971__A1 (.I(_07462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13024__I (.I(_07465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13012__I (.I(_07465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13000__I (.I(_07465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12988__I (.I(_07465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12976__I (.I(_07465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12987__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12985__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12982__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12980__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12978__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12993__A1 (.I(_07470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12991__A1 (.I(_07470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12989__A1 (.I(_07470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12986__A1 (.I(_07470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12984__A1 (.I(_07470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12999__A2 (.I(_07473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12997__A2 (.I(_07473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12994__A2 (.I(_07473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12992__A2 (.I(_07473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12990__A2 (.I(_07473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13005__A1 (.I(_07477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13003__A1 (.I(_07477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13001__A1 (.I(_07477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12998__A1 (.I(_07477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12996__A1 (.I(_07477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13011__A2 (.I(_07480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13009__A2 (.I(_07480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13006__A2 (.I(_07480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13004__A2 (.I(_07480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13002__A2 (.I(_07480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13017__A1 (.I(_07484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13015__A1 (.I(_07484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13013__A1 (.I(_07484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13010__A1 (.I(_07484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13008__A1 (.I(_07484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13023__A2 (.I(_07487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13021__A2 (.I(_07487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13018__A2 (.I(_07487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13016__A2 (.I(_07487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13014__A2 (.I(_07487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13029__A1 (.I(_07491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13027__A1 (.I(_07491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13025__A1 (.I(_07491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13022__A1 (.I(_07491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13020__A1 (.I(_07491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13034__A2 (.I(_07494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13032__A2 (.I(_07494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13030__A2 (.I(_07494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13028__A2 (.I(_07494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13026__A2 (.I(_07494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13397__A1 (.I(_07502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13317__A1 (.I(_07502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13237__A1 (.I(_07502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13157__A1 (.I(_07502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13046__A1 (.I(_07502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13123__I (.I(_07503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13106__I (.I(_07503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13043__I (.I(_07503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13041__I (.I(_07503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13149__A1 (.I(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13146__A1 (.I(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13143__A1 (.I(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13140__A1 (.I(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13042__I (.I(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13059__A2 (.I(_07505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13056__A2 (.I(_07505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13052__A2 (.I(_07505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13049__A2 (.I(_07505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13046__A2 (.I(_07505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13089__I (.I(_07506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13072__I (.I(_07506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13061__I (.I(_07506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13054__I (.I(_07506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13044__I (.I(_07506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13150__A2 (.I(_07507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13147__A2 (.I(_07507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13051__A1 (.I(_07507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13048__A1 (.I(_07507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13045__A1 (.I(_07507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13399__A1 (.I(_07509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13319__A1 (.I(_07509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13239__A1 (.I(_07509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13159__A1 (.I(_07509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13049__A1 (.I(_07509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13401__A1 (.I(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13321__A1 (.I(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13241__A1 (.I(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13161__A1 (.I(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13052__A1 (.I(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13404__A1 (.I(_07513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13324__A1 (.I(_07513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13244__A1 (.I(_07513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13164__A1 (.I(_07513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13056__A1 (.I(_07513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13069__A1 (.I(_07514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13066__A1 (.I(_07514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13063__A1 (.I(_07514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13058__A1 (.I(_07514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13055__A1 (.I(_07514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13406__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13326__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13246__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13166__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13059__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13410__A1 (.I(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13330__A1 (.I(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13250__A1 (.I(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13170__A1 (.I(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A1 (.I(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13130__I (.I(_07519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13113__I (.I(_07519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13096__I (.I(_07519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13079__I (.I(_07519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__I (.I(_07519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13077__A2 (.I(_07520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13074__A2 (.I(_07520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13070__A2 (.I(_07520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13067__A2 (.I(_07520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A2 (.I(_07520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13412__A1 (.I(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13332__A1 (.I(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13252__A1 (.I(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13172__A1 (.I(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13067__A1 (.I(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13414__A1 (.I(_07524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13334__A1 (.I(_07524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13254__A1 (.I(_07524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13174__A1 (.I(_07524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13070__A1 (.I(_07524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13417__A1 (.I(_07526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13337__A1 (.I(_07526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13257__A1 (.I(_07526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13177__A1 (.I(_07526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13074__A1 (.I(_07526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13086__A1 (.I(_07527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13083__A1 (.I(_07527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13080__A1 (.I(_07527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13076__A1 (.I(_07527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13073__A1 (.I(_07527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13419__A1 (.I(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13339__A1 (.I(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13259__A1 (.I(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13179__A1 (.I(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13077__A1 (.I(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__A1 (.I(_07531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13342__A1 (.I(_07531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13262__A1 (.I(_07531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13182__A1 (.I(_07531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13081__A1 (.I(_07531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13094__A2 (.I(_07532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13091__A2 (.I(_07532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__A2 (.I(_07532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13084__A2 (.I(_07532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13081__A2 (.I(_07532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13424__A1 (.I(_07534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13344__A1 (.I(_07534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13264__A1 (.I(_07534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13184__A1 (.I(_07534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13084__A1 (.I(_07534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13426__A1 (.I(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__A1 (.I(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13266__A1 (.I(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13186__A1 (.I(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__A1 (.I(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13429__A1 (.I(_07538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13349__A1 (.I(_07538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13269__A1 (.I(_07538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13189__A1 (.I(_07538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13091__A1 (.I(_07538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13103__A1 (.I(_07539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13100__A1 (.I(_07539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13097__A1 (.I(_07539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13093__A1 (.I(_07539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13090__A1 (.I(_07539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13431__A1 (.I(_07541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13351__A1 (.I(_07541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__A1 (.I(_07541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13191__A1 (.I(_07541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13094__A1 (.I(_07541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13434__A1 (.I(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13354__A1 (.I(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13274__A1 (.I(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13194__A1 (.I(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13098__A1 (.I(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13111__A2 (.I(_07544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13108__A2 (.I(_07544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13104__A2 (.I(_07544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13101__A2 (.I(_07544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13098__A2 (.I(_07544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13436__A1 (.I(_07546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13356__A1 (.I(_07546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13276__A1 (.I(_07546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13196__A1 (.I(_07546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13101__A1 (.I(_07546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13438__A1 (.I(_07548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13358__A1 (.I(_07548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13278__A1 (.I(_07548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13198__A1 (.I(_07548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13104__A1 (.I(_07548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13441__A1 (.I(_07550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13361__A1 (.I(_07550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13281__A1 (.I(_07550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13201__A1 (.I(_07550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13108__A1 (.I(_07550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13120__A1 (.I(_07551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13117__A1 (.I(_07551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13114__A1 (.I(_07551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13110__A1 (.I(_07551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13107__A1 (.I(_07551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13443__A1 (.I(_07553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13363__A1 (.I(_07553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13283__A1 (.I(_07553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__A1 (.I(_07553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13111__A1 (.I(_07553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13446__A1 (.I(_07555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__A1 (.I(_07555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13286__A1 (.I(_07555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13206__A1 (.I(_07555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13115__A1 (.I(_07555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13128__A2 (.I(_07556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13125__A2 (.I(_07556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13121__A2 (.I(_07556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13118__A2 (.I(_07556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13115__A2 (.I(_07556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13448__A1 (.I(_07558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13368__A1 (.I(_07558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13288__A1 (.I(_07558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13208__A1 (.I(_07558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13118__A1 (.I(_07558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13450__A1 (.I(_07560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13370__A1 (.I(_07560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13290__A1 (.I(_07560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13210__A1 (.I(_07560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13121__A1 (.I(_07560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13453__A1 (.I(_07562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13373__A1 (.I(_07562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13293__A1 (.I(_07562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13213__A1 (.I(_07562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13125__A1 (.I(_07562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13137__A1 (.I(_07563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13134__A1 (.I(_07563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13131__A1 (.I(_07563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13127__A1 (.I(_07563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13124__A1 (.I(_07563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13455__A1 (.I(_07565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13375__A1 (.I(_07565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13295__A1 (.I(_07565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13215__A1 (.I(_07565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13128__A1 (.I(_07565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13458__A1 (.I(_07567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13378__A1 (.I(_07567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13298__A1 (.I(_07567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13218__A1 (.I(_07567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13132__A1 (.I(_07567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13144__A2 (.I(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13141__A2 (.I(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13138__A2 (.I(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13135__A2 (.I(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13132__A2 (.I(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13460__A1 (.I(_07570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13380__A1 (.I(_07570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13300__A1 (.I(_07570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13220__A1 (.I(_07570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13135__A1 (.I(_07570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13462__A1 (.I(_07572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13382__A1 (.I(_07572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13302__A1 (.I(_07572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13222__A1 (.I(_07572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13138__A1 (.I(_07572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13464__A1 (.I(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13384__A1 (.I(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13304__A1 (.I(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13224__A1 (.I(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13141__A1 (.I(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13466__A1 (.I(_07576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13386__A1 (.I(_07576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13306__A1 (.I(_07576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13226__A1 (.I(_07576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13144__A1 (.I(_07576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13468__A1 (.I(_07578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13388__A1 (.I(_07578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13308__A1 (.I(_07578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13228__A1 (.I(_07578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13147__A1 (.I(_07578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13470__A1 (.I(_07580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13390__A1 (.I(_07580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13310__A1 (.I(_07580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A1 (.I(_07580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13150__A1 (.I(_07580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13211__I (.I(_07582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13199__I (.I(_07582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13154__I (.I(_07582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13152__I (.I(_07582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13229__A1 (.I(_07583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13227__A1 (.I(_07583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13225__A1 (.I(_07583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13223__A1 (.I(_07583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13153__I (.I(_07583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13166__A2 (.I(_07584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13164__A2 (.I(_07584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13161__A2 (.I(_07584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13159__A2 (.I(_07584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13157__A2 (.I(_07584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13187__I (.I(_07585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13175__I (.I(_07585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13167__I (.I(_07585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13162__I (.I(_07585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13155__I (.I(_07585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A2 (.I(_07586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13228__A2 (.I(_07586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13160__A1 (.I(_07586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13158__A1 (.I(_07586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13156__A1 (.I(_07586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13173__A1 (.I(_07590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13171__A1 (.I(_07590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13169__A1 (.I(_07590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13165__A1 (.I(_07590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13163__A1 (.I(_07590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13216__I (.I(_07593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13204__I (.I(_07593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13192__I (.I(_07593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13180__I (.I(_07593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13168__I (.I(_07593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13179__A2 (.I(_07594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13177__A2 (.I(_07594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13174__A2 (.I(_07594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13172__A2 (.I(_07594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13170__A2 (.I(_07594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13185__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13183__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13181__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13178__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13176__A1 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13191__A2 (.I(_07601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13189__A2 (.I(_07601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13186__A2 (.I(_07601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13184__A2 (.I(_07601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13182__A2 (.I(_07601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13197__A1 (.I(_07605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13195__A1 (.I(_07605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13193__A1 (.I(_07605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13190__A1 (.I(_07605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13188__A1 (.I(_07605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__A2 (.I(_07608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13201__A2 (.I(_07608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13198__A2 (.I(_07608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13196__A2 (.I(_07608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13194__A2 (.I(_07608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13209__A1 (.I(_07612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13207__A1 (.I(_07612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13205__A1 (.I(_07612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13202__A1 (.I(_07612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13200__A1 (.I(_07612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13215__A2 (.I(_07615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13213__A2 (.I(_07615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13210__A2 (.I(_07615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13208__A2 (.I(_07615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13206__A2 (.I(_07615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13221__A1 (.I(_07619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13219__A1 (.I(_07619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13217__A1 (.I(_07619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13214__A1 (.I(_07619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13212__A1 (.I(_07619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13226__A2 (.I(_07622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13224__A2 (.I(_07622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13222__A2 (.I(_07622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13220__A2 (.I(_07622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13218__A2 (.I(_07622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13291__I (.I(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13279__I (.I(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13234__I (.I(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13232__I (.I(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13309__A1 (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13307__A1 (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13305__A1 (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13303__A1 (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13233__I (.I(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13246__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13244__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13241__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13239__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13237__A2 (.I(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13267__I (.I(_07633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13255__I (.I(_07633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13247__I (.I(_07633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13242__I (.I(_07633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13235__I (.I(_07633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13310__A2 (.I(_07634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13308__A2 (.I(_07634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13240__A1 (.I(_07634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13238__A1 (.I(_07634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13236__A1 (.I(_07634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13253__A1 (.I(_07638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13251__A1 (.I(_07638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13249__A1 (.I(_07638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13245__A1 (.I(_07638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13243__A1 (.I(_07638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13296__I (.I(_07641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13284__I (.I(_07641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13272__I (.I(_07641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13260__I (.I(_07641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13248__I (.I(_07641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13259__A2 (.I(_07642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13257__A2 (.I(_07642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13254__A2 (.I(_07642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13252__A2 (.I(_07642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13250__A2 (.I(_07642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13265__A1 (.I(_07646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13263__A1 (.I(_07646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13261__A1 (.I(_07646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13258__A1 (.I(_07646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13256__A1 (.I(_07646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__A2 (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13269__A2 (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13266__A2 (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13264__A2 (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13262__A2 (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13277__A1 (.I(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13275__A1 (.I(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13273__A1 (.I(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13270__A1 (.I(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13268__A1 (.I(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13283__A2 (.I(_07656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13281__A2 (.I(_07656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13278__A2 (.I(_07656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13276__A2 (.I(_07656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13274__A2 (.I(_07656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13289__A1 (.I(_07660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13287__A1 (.I(_07660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13285__A1 (.I(_07660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13282__A1 (.I(_07660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13280__A1 (.I(_07660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13295__A2 (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13293__A2 (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13290__A2 (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13288__A2 (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13286__A2 (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13301__A1 (.I(_07667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13299__A1 (.I(_07667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13297__A1 (.I(_07667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13294__A1 (.I(_07667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13292__A1 (.I(_07667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13306__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13304__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13302__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13300__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13298__A2 (.I(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13371__I (.I(_07678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13359__I (.I(_07678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13314__I (.I(_07678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13312__I (.I(_07678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__A1 (.I(_07679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13387__A1 (.I(_07679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13385__A1 (.I(_07679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13383__A1 (.I(_07679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13313__I (.I(_07679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13326__A2 (.I(_07680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13324__A2 (.I(_07680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13321__A2 (.I(_07680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13319__A2 (.I(_07680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13317__A2 (.I(_07680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13347__I (.I(_07681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13335__I (.I(_07681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13327__I (.I(_07681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13322__I (.I(_07681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13315__I (.I(_07681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13390__A2 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13388__A2 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13320__A1 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13318__A1 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13316__A1 (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13333__A1 (.I(_07686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13331__A1 (.I(_07686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13329__A1 (.I(_07686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13325__A1 (.I(_07686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13323__A1 (.I(_07686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13376__I (.I(_07689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13364__I (.I(_07689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13352__I (.I(_07689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13340__I (.I(_07689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13328__I (.I(_07689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13339__A2 (.I(_07690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13337__A2 (.I(_07690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13334__A2 (.I(_07690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13332__A2 (.I(_07690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13330__A2 (.I(_07690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13345__A1 (.I(_07694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13343__A1 (.I(_07694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13341__A1 (.I(_07694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13338__A1 (.I(_07694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A1 (.I(_07694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13351__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13349__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13344__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13342__A2 (.I(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13357__A1 (.I(_07701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13355__A1 (.I(_07701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13353__A1 (.I(_07701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13350__A1 (.I(_07701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13348__A1 (.I(_07701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13363__A2 (.I(_07704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13361__A2 (.I(_07704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13358__A2 (.I(_07704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13356__A2 (.I(_07704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13354__A2 (.I(_07704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13369__A1 (.I(_07708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13367__A1 (.I(_07708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__A1 (.I(_07708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13362__A1 (.I(_07708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13360__A1 (.I(_07708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13375__A2 (.I(_07711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13373__A2 (.I(_07711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13370__A2 (.I(_07711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13368__A2 (.I(_07711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__A2 (.I(_07711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13381__A1 (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13379__A1 (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__A1 (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13374__A1 (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13372__A1 (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13386__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13384__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13382__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13380__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13378__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13451__I (.I(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13439__I (.I(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13394__I (.I(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13392__I (.I(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13469__A1 (.I(_07727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13467__A1 (.I(_07727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13465__A1 (.I(_07727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13463__A1 (.I(_07727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13393__I (.I(_07727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13406__A2 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13404__A2 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13401__A2 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13399__A2 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13397__A2 (.I(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13427__I (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13415__I (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13407__I (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13402__I (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13395__I (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13470__A2 (.I(_07730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13468__A2 (.I(_07730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13400__A1 (.I(_07730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13398__A1 (.I(_07730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13396__A1 (.I(_07730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13413__A1 (.I(_07734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13411__A1 (.I(_07734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13409__A1 (.I(_07734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13405__A1 (.I(_07734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13403__A1 (.I(_07734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13456__I (.I(_07737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13444__I (.I(_07737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13432__I (.I(_07737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13420__I (.I(_07737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13408__I (.I(_07737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13419__A2 (.I(_07738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13417__A2 (.I(_07738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13414__A2 (.I(_07738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13412__A2 (.I(_07738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13410__A2 (.I(_07738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13425__A1 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13423__A1 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13421__A1 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13418__A1 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13416__A1 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13431__A2 (.I(_07745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13429__A2 (.I(_07745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13426__A2 (.I(_07745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13424__A2 (.I(_07745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__A2 (.I(_07745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13437__A1 (.I(_07749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13435__A1 (.I(_07749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13433__A1 (.I(_07749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13430__A1 (.I(_07749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13428__A1 (.I(_07749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13443__A2 (.I(_07752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13441__A2 (.I(_07752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13438__A2 (.I(_07752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13436__A2 (.I(_07752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13434__A2 (.I(_07752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13449__A1 (.I(_07756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13447__A1 (.I(_07756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13445__A1 (.I(_07756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13442__A1 (.I(_07756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13440__A1 (.I(_07756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13455__A2 (.I(_07759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13453__A2 (.I(_07759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13450__A2 (.I(_07759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13448__A2 (.I(_07759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13446__A2 (.I(_07759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13461__A1 (.I(_07763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13459__A1 (.I(_07763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13457__A1 (.I(_07763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13454__A1 (.I(_07763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13452__A1 (.I(_07763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13466__A2 (.I(_07766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13464__A2 (.I(_07766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13462__A2 (.I(_07766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13460__A2 (.I(_07766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13458__A2 (.I(_07766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(addrD[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(addrD[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(addrD[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(addrD[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(addrD[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(addrS[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(addrS[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(addrS[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(addrS[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(addrS[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(new_value[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(new_value[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(new_value[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(new_value[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(new_value[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(new_value[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(new_value[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(new_value[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(new_value[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(new_value[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(new_value[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(new_value[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(new_value[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(new_value[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(new_value[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(new_value[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(new_value[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(new_value[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(new_value[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(new_value[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(new_value[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(new_value[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(new_value[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(new_value[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(new_value[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(new_value[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(new_value[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(new_value[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(new_value[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(new_value[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(new_value[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(new_value[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14508__A2 (.I(\register_file[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__A2 (.I(\register_file[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A2 (.I(\register_file[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14594__A2 (.I(\register_file[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__A2 (.I(\register_file[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A2 (.I(\register_file[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14679__A2 (.I(\register_file[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__A2 (.I(\register_file[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A2 (.I(\register_file[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14767__A2 (.I(\register_file[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__A2 (.I(\register_file[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(\register_file[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14849__A2 (.I(\register_file[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__A2 (.I(\register_file[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A2 (.I(\register_file[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14930__A2 (.I(\register_file[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11625__A2 (.I(\register_file[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A2 (.I(\register_file[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15101__A2 (.I(\register_file[10][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11629__A2 (.I(\register_file[10][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A2 (.I(\register_file[10][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15187__A2 (.I(\register_file[10][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__A2 (.I(\register_file[10][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A2 (.I(\register_file[10][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15269__A2 (.I(\register_file[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__A2 (.I(\register_file[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A2 (.I(\register_file[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__A2 (.I(\register_file[10][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(\register_file[10][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A2 (.I(\register_file[10][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14345__A2 (.I(\register_file[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__A2 (.I(\register_file[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A2 (.I(\register_file[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14427__A2 (.I(\register_file[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__A2 (.I(\register_file[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(\register_file[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15608__A2 (.I(\register_file[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__A2 (.I(\register_file[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A2 (.I(\register_file[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__A2 (.I(\register_file[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A2 (.I(\register_file[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A2 (.I(\register_file[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__A2 (.I(\register_file[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A2 (.I(\register_file[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A2 (.I(\register_file[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__A2 (.I(\register_file[11][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A2 (.I(\register_file[11][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A2 (.I(\register_file[11][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14168__A2 (.I(\register_file[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A2 (.I(\register_file[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(\register_file[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14511__A2 (.I(\register_file[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A2 (.I(\register_file[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A2 (.I(\register_file[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14598__A2 (.I(\register_file[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A2 (.I(\register_file[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A2 (.I(\register_file[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15526__A2 (.I(\register_file[12][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__A2 (.I(\register_file[12][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A2 (.I(\register_file[12][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A2 (.I(\register_file[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A2 (.I(\register_file[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A2 (.I(\register_file[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14349__A2 (.I(\register_file[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A2 (.I(\register_file[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A2 (.I(\register_file[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14512__A2 (.I(\register_file[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A2 (.I(\register_file[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__A2 (.I(\register_file[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14599__A2 (.I(\register_file[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A2 (.I(\register_file[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A2 (.I(\register_file[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14685__A2 (.I(\register_file[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A2 (.I(\register_file[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(\register_file[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14772__A2 (.I(\register_file[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A2 (.I(\register_file[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A2 (.I(\register_file[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14853__A2 (.I(\register_file[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A2 (.I(\register_file[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A2 (.I(\register_file[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14934__A2 (.I(\register_file[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A2 (.I(\register_file[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A2 (.I(\register_file[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15021__A2 (.I(\register_file[13][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A2 (.I(\register_file[13][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A2 (.I(\register_file[13][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15107__A2 (.I(\register_file[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A2 (.I(\register_file[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__A2 (.I(\register_file[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15192__A2 (.I(\register_file[13][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A2 (.I(\register_file[13][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A2 (.I(\register_file[13][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15273__A2 (.I(\register_file[13][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A2 (.I(\register_file[13][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A2 (.I(\register_file[13][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15354__A2 (.I(\register_file[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A2 (.I(\register_file[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A2 (.I(\register_file[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15442__A2 (.I(\register_file[13][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11207__A2 (.I(\register_file[13][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A2 (.I(\register_file[13][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15529__A2 (.I(\register_file[13][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A2 (.I(\register_file[13][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A2 (.I(\register_file[13][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A2 (.I(\register_file[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A2 (.I(\register_file[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A2 (.I(\register_file[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__A2 (.I(\register_file[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A2 (.I(\register_file[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A2 (.I(\register_file[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A2 (.I(\register_file[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A2 (.I(\register_file[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A2 (.I(\register_file[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A2 (.I(\register_file[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A2 (.I(\register_file[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A2 (.I(\register_file[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A2 (.I(\register_file[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A2 (.I(\register_file[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(\register_file[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13917__A2 (.I(\register_file[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A2 (.I(\register_file[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A2 (.I(\register_file[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14002__A2 (.I(\register_file[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__A2 (.I(\register_file[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A2 (.I(\register_file[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14085__A2 (.I(\register_file[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A2 (.I(\register_file[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(\register_file[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14175__A2 (.I(\register_file[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A2 (.I(\register_file[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(\register_file[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14263__A2 (.I(\register_file[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A2 (.I(\register_file[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A2 (.I(\register_file[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14350__A2 (.I(\register_file[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A2 (.I(\register_file[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A2 (.I(\register_file[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14431__A2 (.I(\register_file[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A2 (.I(\register_file[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A2 (.I(\register_file[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13619__A2 (.I(\register_file[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13236__A2 (.I(\register_file[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A2 (.I(\register_file[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14515__A2 (.I(\register_file[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13261__A2 (.I(\register_file[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A2 (.I(\register_file[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14601__A2 (.I(\register_file[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13263__A2 (.I(\register_file[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A2 (.I(\register_file[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14937__A2 (.I(\register_file[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13273__A2 (.I(\register_file[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A2 (.I(\register_file[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13737__A2 (.I(\register_file[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13238__A2 (.I(\register_file[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A2 (.I(\register_file[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15357__A2 (.I(\register_file[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13285__A2 (.I(\register_file[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A2 (.I(\register_file[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15444__A2 (.I(\register_file[14][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13287__A2 (.I(\register_file[14][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__A2 (.I(\register_file[14][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15531__A2 (.I(\register_file[14][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13289__A2 (.I(\register_file[14][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A2 (.I(\register_file[14][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13292__A2 (.I(\register_file[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A2 (.I(\register_file[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A2 (.I(\register_file[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13294__A2 (.I(\register_file[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A2 (.I(\register_file[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__A2 (.I(\register_file[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13297__A2 (.I(\register_file[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A2 (.I(\register_file[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A2 (.I(\register_file[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13299__A2 (.I(\register_file[14][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A2 (.I(\register_file[14][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(\register_file[14][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13301__A2 (.I(\register_file[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A2 (.I(\register_file[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A2 (.I(\register_file[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13305__A2 (.I(\register_file[14][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A2 (.I(\register_file[14][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A2 (.I(\register_file[14][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13828__A2 (.I(\register_file[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13240__A2 (.I(\register_file[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A2 (.I(\register_file[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13309__A2 (.I(\register_file[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A2 (.I(\register_file[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A2 (.I(\register_file[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13919__A2 (.I(\register_file[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13243__A2 (.I(\register_file[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(\register_file[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14004__A2 (.I(\register_file[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13245__A2 (.I(\register_file[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A2 (.I(\register_file[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14088__A2 (.I(\register_file[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13249__A2 (.I(\register_file[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A2 (.I(\register_file[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14177__A2 (.I(\register_file[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13251__A2 (.I(\register_file[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A2 (.I(\register_file[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14265__A2 (.I(\register_file[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13253__A2 (.I(\register_file[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A2 (.I(\register_file[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14352__A2 (.I(\register_file[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13256__A2 (.I(\register_file[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A2 (.I(\register_file[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14433__A2 (.I(\register_file[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13258__A2 (.I(\register_file[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A2 (.I(\register_file[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13623__A2 (.I(\register_file[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13156__A2 (.I(\register_file[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A2 (.I(\register_file[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14517__A2 (.I(\register_file[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13181__A2 (.I(\register_file[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(\register_file[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14688__A2 (.I(\register_file[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13185__A2 (.I(\register_file[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(\register_file[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13739__A2 (.I(\register_file[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13158__A2 (.I(\register_file[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A2 (.I(\register_file[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15359__A2 (.I(\register_file[15][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13205__A2 (.I(\register_file[15][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A2 (.I(\register_file[15][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15446__A2 (.I(\register_file[15][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13207__A2 (.I(\register_file[15][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A2 (.I(\register_file[15][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15532__A2 (.I(\register_file[15][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13209__A2 (.I(\register_file[15][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A2 (.I(\register_file[15][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13212__A2 (.I(\register_file[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A2 (.I(\register_file[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A2 (.I(\register_file[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13214__A2 (.I(\register_file[15][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A2 (.I(\register_file[15][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A2 (.I(\register_file[15][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13217__A2 (.I(\register_file[15][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A2 (.I(\register_file[15][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A2 (.I(\register_file[15][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13219__A2 (.I(\register_file[15][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A2 (.I(\register_file[15][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A2 (.I(\register_file[15][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13221__A2 (.I(\register_file[15][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__A2 (.I(\register_file[15][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(\register_file[15][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13225__A2 (.I(\register_file[15][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A2 (.I(\register_file[15][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(\register_file[15][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13829__A2 (.I(\register_file[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13160__A2 (.I(\register_file[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A2 (.I(\register_file[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13229__A2 (.I(\register_file[15][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A2 (.I(\register_file[15][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A2 (.I(\register_file[15][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14090__A2 (.I(\register_file[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13169__A2 (.I(\register_file[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A2 (.I(\register_file[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14180__A2 (.I(\register_file[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13171__A2 (.I(\register_file[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A2 (.I(\register_file[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13475__A2 (.I(\register_file[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13045__A2 (.I(\register_file[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(\register_file[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14649__A2 (.I(\register_file[16][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13086__A2 (.I(\register_file[16][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A2 (.I(\register_file[16][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13683__A2 (.I(\register_file[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13048__A2 (.I(\register_file[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A2 (.I(\register_file[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15326__A2 (.I(\register_file[16][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13114__A2 (.I(\register_file[16][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A2 (.I(\register_file[16][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15390__A2 (.I(\register_file[16][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13117__A2 (.I(\register_file[16][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A2 (.I(\register_file[16][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15580__A2 (.I(\register_file[16][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13124__A2 (.I(\register_file[16][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A2 (.I(\register_file[16][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13127__A2 (.I(\register_file[16][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A2 (.I(\register_file[16][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A2 (.I(\register_file[16][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13131__A2 (.I(\register_file[16][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A2 (.I(\register_file[16][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A2 (.I(\register_file[16][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13134__A2 (.I(\register_file[16][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A2 (.I(\register_file[16][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A2 (.I(\register_file[16][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13137__A2 (.I(\register_file[16][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__A2 (.I(\register_file[16][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A2 (.I(\register_file[16][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13140__A2 (.I(\register_file[16][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A2 (.I(\register_file[16][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A2 (.I(\register_file[16][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13143__A2 (.I(\register_file[16][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A2 (.I(\register_file[16][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A2 (.I(\register_file[16][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13769__A2 (.I(\register_file[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13051__A2 (.I(\register_file[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A2 (.I(\register_file[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13146__A2 (.I(\register_file[16][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A2 (.I(\register_file[16][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A2 (.I(\register_file[16][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13149__A2 (.I(\register_file[16][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A2 (.I(\register_file[16][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A2 (.I(\register_file[16][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13859__A2 (.I(\register_file[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13055__A2 (.I(\register_file[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(\register_file[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13968__A2 (.I(\register_file[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13058__A2 (.I(\register_file[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A2 (.I(\register_file[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14057__A2 (.I(\register_file[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13063__A2 (.I(\register_file[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A2 (.I(\register_file[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14140__A2 (.I(\register_file[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13066__A2 (.I(\register_file[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A2 (.I(\register_file[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14226__A2 (.I(\register_file[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13069__A2 (.I(\register_file[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A2 (.I(\register_file[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14315__A2 (.I(\register_file[16][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13073__A2 (.I(\register_file[16][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A2 (.I(\register_file[16][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14399__A2 (.I(\register_file[16][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13076__A2 (.I(\register_file[16][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A2 (.I(\register_file[16][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14485__A2 (.I(\register_file[17][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12989__A2 (.I(\register_file[17][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A2 (.I(\register_file[17][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14567__A2 (.I(\register_file[17][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12991__A2 (.I(\register_file[17][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A2 (.I(\register_file[17][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14651__A2 (.I(\register_file[17][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12993__A2 (.I(\register_file[17][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A2 (.I(\register_file[17][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14738__A2 (.I(\register_file[17][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12996__A2 (.I(\register_file[17][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A2 (.I(\register_file[17][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14822__A2 (.I(\register_file[17][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12998__A2 (.I(\register_file[17][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(\register_file[17][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14907__A2 (.I(\register_file[17][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13001__A2 (.I(\register_file[17][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A2 (.I(\register_file[17][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14989__A2 (.I(\register_file[17][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13003__A2 (.I(\register_file[17][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A2 (.I(\register_file[17][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15073__A2 (.I(\register_file[17][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13005__A2 (.I(\register_file[17][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A2 (.I(\register_file[17][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15139__A2 (.I(\register_file[17][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13008__A2 (.I(\register_file[17][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A2 (.I(\register_file[17][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15222__A2 (.I(\register_file[17][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13010__A2 (.I(\register_file[17][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A2 (.I(\register_file[17][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15327__A2 (.I(\register_file[17][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13013__A2 (.I(\register_file[17][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A2 (.I(\register_file[17][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15391__A2 (.I(\register_file[17][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13015__A2 (.I(\register_file[17][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__A2 (.I(\register_file[17][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15476__A2 (.I(\register_file[17][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13017__A2 (.I(\register_file[17][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A2 (.I(\register_file[17][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15581__A2 (.I(\register_file[17][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13020__A2 (.I(\register_file[17][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A2 (.I(\register_file[17][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13022__A2 (.I(\register_file[17][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A2 (.I(\register_file[17][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A2 (.I(\register_file[17][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13031__A2 (.I(\register_file[17][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A2 (.I(\register_file[17][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A2 (.I(\register_file[17][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13035__A2 (.I(\register_file[17][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A2 (.I(\register_file[17][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A2 (.I(\register_file[17][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13860__A2 (.I(\register_file[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12971__A2 (.I(\register_file[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(\register_file[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13969__A2 (.I(\register_file[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12973__A2 (.I(\register_file[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A2 (.I(\register_file[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14058__A2 (.I(\register_file[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12977__A2 (.I(\register_file[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A2 (.I(\register_file[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14141__A2 (.I(\register_file[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12979__A2 (.I(\register_file[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A2 (.I(\register_file[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14228__A2 (.I(\register_file[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12981__A2 (.I(\register_file[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A2 (.I(\register_file[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14316__A2 (.I(\register_file[17][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12984__A2 (.I(\register_file[17][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(\register_file[17][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14400__A2 (.I(\register_file[17][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12986__A2 (.I(\register_file[17][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A2 (.I(\register_file[17][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14490__A2 (.I(\register_file[18][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__A2 (.I(\register_file[18][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A2 (.I(\register_file[18][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14572__A2 (.I(\register_file[18][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12911__A2 (.I(\register_file[18][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__A2 (.I(\register_file[18][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14657__A2 (.I(\register_file[18][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12913__A2 (.I(\register_file[18][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A2 (.I(\register_file[18][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14745__A2 (.I(\register_file[18][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__A2 (.I(\register_file[18][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A2 (.I(\register_file[18][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14828__A2 (.I(\register_file[18][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12918__A2 (.I(\register_file[18][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(\register_file[18][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14912__A2 (.I(\register_file[18][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12921__A2 (.I(\register_file[18][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A2 (.I(\register_file[18][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14994__A2 (.I(\register_file[18][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12923__A2 (.I(\register_file[18][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A2 (.I(\register_file[18][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15079__A2 (.I(\register_file[18][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12925__A2 (.I(\register_file[18][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A2 (.I(\register_file[18][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15145__A2 (.I(\register_file[18][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12928__A2 (.I(\register_file[18][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A2 (.I(\register_file[18][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15227__A2 (.I(\register_file[18][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12930__A2 (.I(\register_file[18][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A2 (.I(\register_file[18][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15332__A2 (.I(\register_file[18][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12933__A2 (.I(\register_file[18][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A2 (.I(\register_file[18][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15396__A2 (.I(\register_file[18][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12935__A2 (.I(\register_file[18][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A2 (.I(\register_file[18][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15482__A2 (.I(\register_file[18][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12937__A2 (.I(\register_file[18][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__A2 (.I(\register_file[18][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15587__A2 (.I(\register_file[18][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12940__A2 (.I(\register_file[18][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A2 (.I(\register_file[18][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12942__A2 (.I(\register_file[18][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A2 (.I(\register_file[18][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A2 (.I(\register_file[18][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12945__A2 (.I(\register_file[18][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A2 (.I(\register_file[18][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A2 (.I(\register_file[18][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__A2 (.I(\register_file[18][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A2 (.I(\register_file[18][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A2 (.I(\register_file[18][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12953__A2 (.I(\register_file[18][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A2 (.I(\register_file[18][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A2 (.I(\register_file[18][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12957__A2 (.I(\register_file[18][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__A2 (.I(\register_file[18][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A2 (.I(\register_file[18][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13866__A2 (.I(\register_file[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12891__A2 (.I(\register_file[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A2 (.I(\register_file[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13976__A2 (.I(\register_file[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12893__A2 (.I(\register_file[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A2 (.I(\register_file[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14063__A2 (.I(\register_file[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12897__A2 (.I(\register_file[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A2 (.I(\register_file[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14146__A2 (.I(\register_file[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12899__A2 (.I(\register_file[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A2 (.I(\register_file[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14234__A2 (.I(\register_file[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12901__A2 (.I(\register_file[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A2 (.I(\register_file[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14323__A2 (.I(\register_file[18][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12904__A2 (.I(\register_file[18][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(\register_file[18][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14406__A2 (.I(\register_file[18][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12906__A2 (.I(\register_file[18][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A2 (.I(\register_file[18][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14656__A2 (.I(\register_file[19][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__A2 (.I(\register_file[19][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(\register_file[19][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14993__A2 (.I(\register_file[19][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__A2 (.I(\register_file[19][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A2 (.I(\register_file[19][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15226__A2 (.I(\register_file[19][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A2 (.I(\register_file[19][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A2 (.I(\register_file[19][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15395__A2 (.I(\register_file[19][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A2 (.I(\register_file[19][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A2 (.I(\register_file[19][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15585__A2 (.I(\register_file[19][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A2 (.I(\register_file[19][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__A2 (.I(\register_file[19][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__A2 (.I(\register_file[19][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A2 (.I(\register_file[19][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A2 (.I(\register_file[19][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__A2 (.I(\register_file[19][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A2 (.I(\register_file[19][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(\register_file[19][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A2 (.I(\register_file[19][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A2 (.I(\register_file[19][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A2 (.I(\register_file[19][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A2 (.I(\register_file[19][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A2 (.I(\register_file[19][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__A2 (.I(\register_file[19][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A2 (.I(\register_file[19][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__A2 (.I(\register_file[19][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A2 (.I(\register_file[19][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13865__A2 (.I(\register_file[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A2 (.I(\register_file[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(\register_file[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13975__A2 (.I(\register_file[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A2 (.I(\register_file[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A2 (.I(\register_file[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14233__A2 (.I(\register_file[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A2 (.I(\register_file[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A2 (.I(\register_file[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14405__A2 (.I(\register_file[19][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A2 (.I(\register_file[19][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(\register_file[19][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14539__A2 (.I(\register_file[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12829__A2 (.I(\register_file[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A2 (.I(\register_file[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14626__A2 (.I(\register_file[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12831__A2 (.I(\register_file[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A2 (.I(\register_file[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14710__A2 (.I(\register_file[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12833__A2 (.I(\register_file[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(\register_file[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14795__A2 (.I(\register_file[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12836__A2 (.I(\register_file[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A2 (.I(\register_file[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14877__A2 (.I(\register_file[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12838__A2 (.I(\register_file[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A2 (.I(\register_file[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14961__A2 (.I(\register_file[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12841__A2 (.I(\register_file[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(\register_file[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15048__A2 (.I(\register_file[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12843__A2 (.I(\register_file[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(\register_file[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15132__A2 (.I(\register_file[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__A2 (.I(\register_file[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A2 (.I(\register_file[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15215__A2 (.I(\register_file[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12848__A2 (.I(\register_file[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A2 (.I(\register_file[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15297__A2 (.I(\register_file[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12850__A2 (.I(\register_file[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A2 (.I(\register_file[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13763__A2 (.I(\register_file[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12806__A2 (.I(\register_file[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A2 (.I(\register_file[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15381__A2 (.I(\register_file[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12853__A2 (.I(\register_file[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A2 (.I(\register_file[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15469__A2 (.I(\register_file[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12855__A2 (.I(\register_file[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__A2 (.I(\register_file[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15554__A2 (.I(\register_file[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12857__A2 (.I(\register_file[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A2 (.I(\register_file[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12860__A2 (.I(\register_file[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A2 (.I(\register_file[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A2 (.I(\register_file[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12862__A2 (.I(\register_file[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A2 (.I(\register_file[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A2 (.I(\register_file[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12865__A2 (.I(\register_file[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A2 (.I(\register_file[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A2 (.I(\register_file[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12867__A2 (.I(\register_file[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A2 (.I(\register_file[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A2 (.I(\register_file[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__A2 (.I(\register_file[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__A2 (.I(\register_file[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A2 (.I(\register_file[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12875__A2 (.I(\register_file[1][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A2 (.I(\register_file[1][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__A2 (.I(\register_file[1][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14112__A2 (.I(\register_file[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12817__A2 (.I(\register_file[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A2 (.I(\register_file[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14203__A2 (.I(\register_file[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12819__A2 (.I(\register_file[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A2 (.I(\register_file[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14288__A2 (.I(\register_file[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12821__A2 (.I(\register_file[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A2 (.I(\register_file[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14373__A2 (.I(\register_file[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12824__A2 (.I(\register_file[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A2 (.I(\register_file[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14455__A2 (.I(\register_file[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12826__A2 (.I(\register_file[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A2 (.I(\register_file[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14493__A2 (.I(\register_file[20][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__A2 (.I(\register_file[20][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A2 (.I(\register_file[20][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14575__A2 (.I(\register_file[20][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12751__A2 (.I(\register_file[20][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A2 (.I(\register_file[20][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14661__A2 (.I(\register_file[20][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12753__A2 (.I(\register_file[20][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A2 (.I(\register_file[20][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14832__A2 (.I(\register_file[20][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12758__A2 (.I(\register_file[20][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A2 (.I(\register_file[20][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14915__A2 (.I(\register_file[20][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12761__A2 (.I(\register_file[20][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(\register_file[20][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14997__A2 (.I(\register_file[20][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12763__A2 (.I(\register_file[20][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A2 (.I(\register_file[20][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15083__A2 (.I(\register_file[20][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12765__A2 (.I(\register_file[20][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A2 (.I(\register_file[20][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15149__A2 (.I(\register_file[20][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12768__A2 (.I(\register_file[20][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A2 (.I(\register_file[20][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15230__A2 (.I(\register_file[20][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12770__A2 (.I(\register_file[20][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__A2 (.I(\register_file[20][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15335__A2 (.I(\register_file[20][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12773__A2 (.I(\register_file[20][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A2 (.I(\register_file[20][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15399__A2 (.I(\register_file[20][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12775__A2 (.I(\register_file[20][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__A2 (.I(\register_file[20][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15485__A2 (.I(\register_file[20][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12777__A2 (.I(\register_file[20][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A2 (.I(\register_file[20][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15590__A2 (.I(\register_file[20][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12780__A2 (.I(\register_file[20][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A2 (.I(\register_file[20][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12782__A2 (.I(\register_file[20][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A2 (.I(\register_file[20][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__A2 (.I(\register_file[20][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12793__A2 (.I(\register_file[20][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A2 (.I(\register_file[20][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A2 (.I(\register_file[20][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13870__A2 (.I(\register_file[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12731__A2 (.I(\register_file[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A2 (.I(\register_file[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13980__A2 (.I(\register_file[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12733__A2 (.I(\register_file[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A2 (.I(\register_file[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14066__A2 (.I(\register_file[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12737__A2 (.I(\register_file[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A2 (.I(\register_file[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14149__A2 (.I(\register_file[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12739__A2 (.I(\register_file[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(\register_file[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14238__A2 (.I(\register_file[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12741__A2 (.I(\register_file[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A2 (.I(\register_file[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14326__A2 (.I(\register_file[20][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12744__A2 (.I(\register_file[20][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A2 (.I(\register_file[20][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14410__A2 (.I(\register_file[20][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12746__A2 (.I(\register_file[20][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A2 (.I(\register_file[20][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14494__A2 (.I(\register_file[21][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12648__A2 (.I(\register_file[21][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A2 (.I(\register_file[21][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14576__A2 (.I(\register_file[21][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12651__A2 (.I(\register_file[21][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A2 (.I(\register_file[21][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14662__A2 (.I(\register_file[21][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12654__A2 (.I(\register_file[21][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A2 (.I(\register_file[21][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14751__A2 (.I(\register_file[21][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12658__A2 (.I(\register_file[21][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A2 (.I(\register_file[21][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14833__A2 (.I(\register_file[21][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__A2 (.I(\register_file[21][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A2 (.I(\register_file[21][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14916__A2 (.I(\register_file[21][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12665__A2 (.I(\register_file[21][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A2 (.I(\register_file[21][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14998__A2 (.I(\register_file[21][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12668__A2 (.I(\register_file[21][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A2 (.I(\register_file[21][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15084__A2 (.I(\register_file[21][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12671__A2 (.I(\register_file[21][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__A2 (.I(\register_file[21][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15150__A2 (.I(\register_file[21][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12675__A2 (.I(\register_file[21][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A2 (.I(\register_file[21][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15232__A2 (.I(\register_file[21][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12678__A2 (.I(\register_file[21][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A2 (.I(\register_file[21][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15336__A2 (.I(\register_file[21][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12682__A2 (.I(\register_file[21][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A2 (.I(\register_file[21][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15400__A2 (.I(\register_file[21][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12685__A2 (.I(\register_file[21][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A2 (.I(\register_file[21][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15486__A2 (.I(\register_file[21][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12688__A2 (.I(\register_file[21][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A2 (.I(\register_file[21][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15593__A2 (.I(\register_file[21][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12692__A2 (.I(\register_file[21][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A2 (.I(\register_file[21][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12714__A2 (.I(\register_file[21][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__A2 (.I(\register_file[21][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__A2 (.I(\register_file[21][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13871__A2 (.I(\register_file[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__A2 (.I(\register_file[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A2 (.I(\register_file[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13981__A2 (.I(\register_file[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__A2 (.I(\register_file[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A2 (.I(\register_file[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14067__A2 (.I(\register_file[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12631__A2 (.I(\register_file[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A2 (.I(\register_file[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14150__A2 (.I(\register_file[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12634__A2 (.I(\register_file[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(\register_file[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14239__A2 (.I(\register_file[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__A2 (.I(\register_file[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(\register_file[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14329__A2 (.I(\register_file[21][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12641__A2 (.I(\register_file[21][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A2 (.I(\register_file[21][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14411__A2 (.I(\register_file[21][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12644__A2 (.I(\register_file[21][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A2 (.I(\register_file[21][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13523__A2 (.I(\register_file[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12532__A2 (.I(\register_file[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A2 (.I(\register_file[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14496__A2 (.I(\register_file[22][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12557__A2 (.I(\register_file[22][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A2 (.I(\register_file[22][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14578__A2 (.I(\register_file[22][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12559__A2 (.I(\register_file[22][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(\register_file[22][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14665__A2 (.I(\register_file[22][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12561__A2 (.I(\register_file[22][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A2 (.I(\register_file[22][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14753__A2 (.I(\register_file[22][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12564__A2 (.I(\register_file[22][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A2 (.I(\register_file[22][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14835__A2 (.I(\register_file[22][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12566__A2 (.I(\register_file[22][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(\register_file[22][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14918__A2 (.I(\register_file[22][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12569__A2 (.I(\register_file[22][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A2 (.I(\register_file[22][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15000__A2 (.I(\register_file[22][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12571__A2 (.I(\register_file[22][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A2 (.I(\register_file[22][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15087__A2 (.I(\register_file[22][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12573__A2 (.I(\register_file[22][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A2 (.I(\register_file[22][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15152__A2 (.I(\register_file[22][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12576__A2 (.I(\register_file[22][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A2 (.I(\register_file[22][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15235__A2 (.I(\register_file[22][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12578__A2 (.I(\register_file[22][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A2 (.I(\register_file[22][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13695__A2 (.I(\register_file[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__A2 (.I(\register_file[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__A2 (.I(\register_file[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15338__A2 (.I(\register_file[22][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12581__A2 (.I(\register_file[22][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A2 (.I(\register_file[22][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15402__A2 (.I(\register_file[22][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__A2 (.I(\register_file[22][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__A2 (.I(\register_file[22][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15488__A2 (.I(\register_file[22][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12585__A2 (.I(\register_file[22][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A2 (.I(\register_file[22][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12599__A2 (.I(\register_file[22][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__A2 (.I(\register_file[22][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A2 (.I(\register_file[22][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13782__A2 (.I(\register_file[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__A2 (.I(\register_file[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A2 (.I(\register_file[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__A2 (.I(\register_file[22][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A2 (.I(\register_file[22][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__A2 (.I(\register_file[22][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12605__A2 (.I(\register_file[22][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A2 (.I(\register_file[22][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A2 (.I(\register_file[22][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14069__A2 (.I(\register_file[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12545__A2 (.I(\register_file[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A2 (.I(\register_file[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14152__A2 (.I(\register_file[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__A2 (.I(\register_file[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A2 (.I(\register_file[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14331__A2 (.I(\register_file[22][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12552__A2 (.I(\register_file[22][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A2 (.I(\register_file[22][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14413__A2 (.I(\register_file[22][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12554__A2 (.I(\register_file[22][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(\register_file[22][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13528__A2 (.I(\register_file[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12452__A2 (.I(\register_file[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A2 (.I(\register_file[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14497__A2 (.I(\register_file[23][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12477__A2 (.I(\register_file[23][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A2 (.I(\register_file[23][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14579__A2 (.I(\register_file[23][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12479__A2 (.I(\register_file[23][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A2 (.I(\register_file[23][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14668__A2 (.I(\register_file[23][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__A2 (.I(\register_file[23][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(\register_file[23][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14754__A2 (.I(\register_file[23][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12484__A2 (.I(\register_file[23][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A2 (.I(\register_file[23][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14836__A2 (.I(\register_file[23][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12486__A2 (.I(\register_file[23][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A2 (.I(\register_file[23][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14919__A2 (.I(\register_file[23][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__A2 (.I(\register_file[23][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(\register_file[23][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15001__A2 (.I(\register_file[23][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12491__A2 (.I(\register_file[23][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A2 (.I(\register_file[23][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15090__A2 (.I(\register_file[23][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12493__A2 (.I(\register_file[23][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A2 (.I(\register_file[23][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15153__A2 (.I(\register_file[23][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12496__A2 (.I(\register_file[23][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A2 (.I(\register_file[23][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15237__A2 (.I(\register_file[23][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12498__A2 (.I(\register_file[23][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A2 (.I(\register_file[23][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13697__A2 (.I(\register_file[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12454__A2 (.I(\register_file[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A2 (.I(\register_file[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15339__A2 (.I(\register_file[23][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12501__A2 (.I(\register_file[23][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__A2 (.I(\register_file[23][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15404__A2 (.I(\register_file[23][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12503__A2 (.I(\register_file[23][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A2 (.I(\register_file[23][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15489__A2 (.I(\register_file[23][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12505__A2 (.I(\register_file[23][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A2 (.I(\register_file[23][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15596__A2 (.I(\register_file[23][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12508__A2 (.I(\register_file[23][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A2 (.I(\register_file[23][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12510__A2 (.I(\register_file[23][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A2 (.I(\register_file[23][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A2 (.I(\register_file[23][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12513__A2 (.I(\register_file[23][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A2 (.I(\register_file[23][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A2 (.I(\register_file[23][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12515__A2 (.I(\register_file[23][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A2 (.I(\register_file[23][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A2 (.I(\register_file[23][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__A2 (.I(\register_file[23][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A2 (.I(\register_file[23][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A2 (.I(\register_file[23][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12519__A2 (.I(\register_file[23][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A2 (.I(\register_file[23][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A2 (.I(\register_file[23][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12521__A2 (.I(\register_file[23][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A2 (.I(\register_file[23][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A2 (.I(\register_file[23][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13783__A2 (.I(\register_file[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12456__A2 (.I(\register_file[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A2 (.I(\register_file[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12523__A2 (.I(\register_file[23][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A2 (.I(\register_file[23][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A2 (.I(\register_file[23][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__A2 (.I(\register_file[23][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__A2 (.I(\register_file[23][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__I (.I(\register_file[23][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13874__A2 (.I(\register_file[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12459__A2 (.I(\register_file[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A2 (.I(\register_file[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13984__A2 (.I(\register_file[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__A2 (.I(\register_file[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A2 (.I(\register_file[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14070__A2 (.I(\register_file[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12465__A2 (.I(\register_file[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A2 (.I(\register_file[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14153__A2 (.I(\register_file[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12467__A2 (.I(\register_file[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A2 (.I(\register_file[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13536__A2 (.I(\register_file[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12372__A2 (.I(\register_file[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A2 (.I(\register_file[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14461__A2 (.I(\register_file[24][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12397__A2 (.I(\register_file[24][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A2 (.I(\register_file[24][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14548__A2 (.I(\register_file[24][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12399__A2 (.I(\register_file[24][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A2 (.I(\register_file[24][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14632__A2 (.I(\register_file[24][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12401__A2 (.I(\register_file[24][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A2 (.I(\register_file[24][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14716__A2 (.I(\register_file[24][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12404__A2 (.I(\register_file[24][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A2 (.I(\register_file[24][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14801__A2 (.I(\register_file[24][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12406__A2 (.I(\register_file[24][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A2 (.I(\register_file[24][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14883__A2 (.I(\register_file[24][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12409__A2 (.I(\register_file[24][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A2 (.I(\register_file[24][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14970__A2 (.I(\register_file[24][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12411__A2 (.I(\register_file[24][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A2 (.I(\register_file[24][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15054__A2 (.I(\register_file[24][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12413__A2 (.I(\register_file[24][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A2 (.I(\register_file[24][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15158__A2 (.I(\register_file[24][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12416__A2 (.I(\register_file[24][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A2 (.I(\register_file[24][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15241__A2 (.I(\register_file[24][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12418__A2 (.I(\register_file[24][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A2 (.I(\register_file[24][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13701__A2 (.I(\register_file[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12374__A2 (.I(\register_file[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A2 (.I(\register_file[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15303__A2 (.I(\register_file[24][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12421__A2 (.I(\register_file[24][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A2 (.I(\register_file[24][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15408__A2 (.I(\register_file[24][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12423__A2 (.I(\register_file[24][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A2 (.I(\register_file[24][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15493__A2 (.I(\register_file[24][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12425__A2 (.I(\register_file[24][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A2 (.I(\register_file[24][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15560__A2 (.I(\register_file[24][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12428__A2 (.I(\register_file[24][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A2 (.I(\register_file[24][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12430__A2 (.I(\register_file[24][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A2 (.I(\register_file[24][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A2 (.I(\register_file[24][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12435__A2 (.I(\register_file[24][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A2 (.I(\register_file[24][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(\register_file[24][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12437__A2 (.I(\register_file[24][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A2 (.I(\register_file[24][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A2 (.I(\register_file[24][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12439__A2 (.I(\register_file[24][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A2 (.I(\register_file[24][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A2 (.I(\register_file[24][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12441__A2 (.I(\register_file[24][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A2 (.I(\register_file[24][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__A2 (.I(\register_file[24][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__A2 (.I(\register_file[24][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A2 (.I(\register_file[24][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A2 (.I(\register_file[24][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12445__A2 (.I(\register_file[24][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__A2 (.I(\register_file[24][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A2 (.I(\register_file[24][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13880__A2 (.I(\register_file[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12379__A2 (.I(\register_file[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A2 (.I(\register_file[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14033__A2 (.I(\register_file[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12385__A2 (.I(\register_file[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A2 (.I(\register_file[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14121__A2 (.I(\register_file[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12387__A2 (.I(\register_file[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(\register_file[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14209__A2 (.I(\register_file[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12389__A2 (.I(\register_file[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A2 (.I(\register_file[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14294__A2 (.I(\register_file[24][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12392__A2 (.I(\register_file[24][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A2 (.I(\register_file[24][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14379__A2 (.I(\register_file[24][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12394__A2 (.I(\register_file[24][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A2 (.I(\register_file[24][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14463__A2 (.I(\register_file[25][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12317__A2 (.I(\register_file[25][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A2 (.I(\register_file[25][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14549__A2 (.I(\register_file[25][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12319__A2 (.I(\register_file[25][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A2 (.I(\register_file[25][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14633__A2 (.I(\register_file[25][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12321__A2 (.I(\register_file[25][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A2 (.I(\register_file[25][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14717__A2 (.I(\register_file[25][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12324__A2 (.I(\register_file[25][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A2 (.I(\register_file[25][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14802__A2 (.I(\register_file[25][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12326__A2 (.I(\register_file[25][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A2 (.I(\register_file[25][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14885__A2 (.I(\register_file[25][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12329__A2 (.I(\register_file[25][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A2 (.I(\register_file[25][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14971__A2 (.I(\register_file[25][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12331__A2 (.I(\register_file[25][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A2 (.I(\register_file[25][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15055__A2 (.I(\register_file[25][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12333__A2 (.I(\register_file[25][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(\register_file[25][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15159__A2 (.I(\register_file[25][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12336__A2 (.I(\register_file[25][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A2 (.I(\register_file[25][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15242__A2 (.I(\register_file[25][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12338__A2 (.I(\register_file[25][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A2 (.I(\register_file[25][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15305__A2 (.I(\register_file[25][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12341__A2 (.I(\register_file[25][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__A2 (.I(\register_file[25][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15409__A2 (.I(\register_file[25][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12343__A2 (.I(\register_file[25][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A2 (.I(\register_file[25][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15495__A2 (.I(\register_file[25][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12345__A2 (.I(\register_file[25][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A2 (.I(\register_file[25][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15561__A2 (.I(\register_file[25][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12348__A2 (.I(\register_file[25][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A2 (.I(\register_file[25][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12350__A2 (.I(\register_file[25][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A2 (.I(\register_file[25][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A2 (.I(\register_file[25][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12355__A2 (.I(\register_file[25][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A2 (.I(\register_file[25][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(\register_file[25][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12357__A2 (.I(\register_file[25][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__A2 (.I(\register_file[25][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A2 (.I(\register_file[25][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12359__A2 (.I(\register_file[25][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A2 (.I(\register_file[25][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(\register_file[25][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12361__A2 (.I(\register_file[25][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A2 (.I(\register_file[25][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A2 (.I(\register_file[25][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12363__A2 (.I(\register_file[25][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A2 (.I(\register_file[25][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A2 (.I(\register_file[25][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__A2 (.I(\register_file[25][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A2 (.I(\register_file[25][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__I (.I(\register_file[25][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13881__A2 (.I(\register_file[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12299__A2 (.I(\register_file[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A2 (.I(\register_file[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14035__A2 (.I(\register_file[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12305__A2 (.I(\register_file[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A2 (.I(\register_file[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14122__A2 (.I(\register_file[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12307__A2 (.I(\register_file[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A2 (.I(\register_file[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14295__A2 (.I(\register_file[25][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12312__A2 (.I(\register_file[25][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A2 (.I(\register_file[25][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14380__A2 (.I(\register_file[25][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12314__A2 (.I(\register_file[25][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A2 (.I(\register_file[25][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13552__A2 (.I(\register_file[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A2 (.I(\register_file[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A2 (.I(\register_file[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14807__A2 (.I(\register_file[26][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A2 (.I(\register_file[26][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A2 (.I(\register_file[26][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13708__A2 (.I(\register_file[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A2 (.I(\register_file[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A2 (.I(\register_file[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15567__A2 (.I(\register_file[26][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A2 (.I(\register_file[26][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A2 (.I(\register_file[26][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__A2 (.I(\register_file[26][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A2 (.I(\register_file[26][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A2 (.I(\register_file[26][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A2 (.I(\register_file[26][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A2 (.I(\register_file[26][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A2 (.I(\register_file[26][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A2 (.I(\register_file[26][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A2 (.I(\register_file[26][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A2 (.I(\register_file[26][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A2 (.I(\register_file[26][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__A2 (.I(\register_file[26][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A2 (.I(\register_file[26][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A2 (.I(\register_file[26][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A2 (.I(\register_file[26][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A2 (.I(\register_file[26][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13796__A2 (.I(\register_file[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A2 (.I(\register_file[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(\register_file[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13888__A2 (.I(\register_file[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__A2 (.I(\register_file[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A2 (.I(\register_file[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14468__A2 (.I(\register_file[27][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A2 (.I(\register_file[27][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A2 (.I(\register_file[27][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14553__A2 (.I(\register_file[27][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__A2 (.I(\register_file[27][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A2 (.I(\register_file[27][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14637__A2 (.I(\register_file[27][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A2 (.I(\register_file[27][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A2 (.I(\register_file[27][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14723__A2 (.I(\register_file[27][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A2 (.I(\register_file[27][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A2 (.I(\register_file[27][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14806__A2 (.I(\register_file[27][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A2 (.I(\register_file[27][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A2 (.I(\register_file[27][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14890__A2 (.I(\register_file[27][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__A2 (.I(\register_file[27][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A2 (.I(\register_file[27][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14975__A2 (.I(\register_file[27][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A2 (.I(\register_file[27][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A2 (.I(\register_file[27][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15059__A2 (.I(\register_file[27][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A2 (.I(\register_file[27][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A2 (.I(\register_file[27][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15163__A2 (.I(\register_file[27][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__A2 (.I(\register_file[27][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A2 (.I(\register_file[27][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15247__A2 (.I(\register_file[27][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A2 (.I(\register_file[27][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A2 (.I(\register_file[27][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15310__A2 (.I(\register_file[27][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A2 (.I(\register_file[27][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A2 (.I(\register_file[27][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15414__A2 (.I(\register_file[27][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__A2 (.I(\register_file[27][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A2 (.I(\register_file[27][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15500__A2 (.I(\register_file[27][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A2 (.I(\register_file[27][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A2 (.I(\register_file[27][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15566__A2 (.I(\register_file[27][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A2 (.I(\register_file[27][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(\register_file[27][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A2 (.I(\register_file[27][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A2 (.I(\register_file[27][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A2 (.I(\register_file[27][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__A2 (.I(\register_file[27][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A2 (.I(\register_file[27][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A2 (.I(\register_file[27][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A2 (.I(\register_file[27][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A2 (.I(\register_file[27][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A2 (.I(\register_file[27][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A2 (.I(\register_file[27][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A2 (.I(\register_file[27][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A2 (.I(\register_file[27][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A2 (.I(\register_file[27][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(\register_file[27][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__A2 (.I(\register_file[27][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13885__A2 (.I(\register_file[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A2 (.I(\register_file[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A2 (.I(\register_file[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13953__A2 (.I(\register_file[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A2 (.I(\register_file[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__A2 (.I(\register_file[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14040__A2 (.I(\register_file[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A2 (.I(\register_file[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A2 (.I(\register_file[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14126__A2 (.I(\register_file[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__A2 (.I(\register_file[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A2 (.I(\register_file[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14214__A2 (.I(\register_file[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A2 (.I(\register_file[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A2 (.I(\register_file[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14301__A2 (.I(\register_file[27][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__A2 (.I(\register_file[27][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A2 (.I(\register_file[27][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14384__A2 (.I(\register_file[27][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A2 (.I(\register_file[27][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A2 (.I(\register_file[27][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14474__A2 (.I(\register_file[28][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A2 (.I(\register_file[28][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A2 (.I(\register_file[28][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14557__A2 (.I(\register_file[28][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(\register_file[28][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A2 (.I(\register_file[28][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14641__A2 (.I(\register_file[28][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A2 (.I(\register_file[28][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A2 (.I(\register_file[28][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14810__A2 (.I(\register_file[28][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A2 (.I(\register_file[28][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A2 (.I(\register_file[28][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14896__A2 (.I(\register_file[28][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A2 (.I(\register_file[28][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A2 (.I(\register_file[28][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15063__A2 (.I(\register_file[28][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__A2 (.I(\register_file[28][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A2 (.I(\register_file[28][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15316__A2 (.I(\register_file[28][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A2 (.I(\register_file[28][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A2 (.I(\register_file[28][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15418__A2 (.I(\register_file[28][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A2 (.I(\register_file[28][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A2 (.I(\register_file[28][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15505__A2 (.I(\register_file[28][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A2 (.I(\register_file[28][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A2 (.I(\register_file[28][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15571__A2 (.I(\register_file[28][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__A2 (.I(\register_file[28][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A2 (.I(\register_file[28][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A2 (.I(\register_file[28][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A2 (.I(\register_file[28][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(\register_file[28][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A2 (.I(\register_file[28][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A2 (.I(\register_file[28][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A2 (.I(\register_file[28][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A2 (.I(\register_file[28][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A2 (.I(\register_file[28][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(\register_file[28][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A2 (.I(\register_file[28][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A2 (.I(\register_file[28][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A2 (.I(\register_file[28][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A2 (.I(\register_file[28][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A2 (.I(\register_file[28][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(\register_file[28][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13891__A2 (.I(\register_file[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A2 (.I(\register_file[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A2 (.I(\register_file[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13957__A2 (.I(\register_file[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A2 (.I(\register_file[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A2 (.I(\register_file[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14047__A2 (.I(\register_file[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__A2 (.I(\register_file[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A2 (.I(\register_file[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14130__A2 (.I(\register_file[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A2 (.I(\register_file[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A2 (.I(\register_file[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14218__A2 (.I(\register_file[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A2 (.I(\register_file[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(\register_file[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14306__A2 (.I(\register_file[28][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A2 (.I(\register_file[28][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A2 (.I(\register_file[28][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14388__A2 (.I(\register_file[28][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A2 (.I(\register_file[28][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A2 (.I(\register_file[28][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13566__A2 (.I(\register_file[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13316__A2 (.I(\register_file[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A2 (.I(\register_file[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14476__A2 (.I(\register_file[29][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13341__A2 (.I(\register_file[29][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A2 (.I(\register_file[29][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14558__A2 (.I(\register_file[29][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13343__A2 (.I(\register_file[29][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A2 (.I(\register_file[29][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14812__A2 (.I(\register_file[29][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13350__A2 (.I(\register_file[29][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__A2 (.I(\register_file[29][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13712__A2 (.I(\register_file[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13318__A2 (.I(\register_file[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A2 (.I(\register_file[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15318__A2 (.I(\register_file[29][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__A2 (.I(\register_file[29][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__A2 (.I(\register_file[29][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15419__A2 (.I(\register_file[29][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13367__A2 (.I(\register_file[29][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A2 (.I(\register_file[29][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15506__A2 (.I(\register_file[29][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13369__A2 (.I(\register_file[29][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A2 (.I(\register_file[29][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15572__A2 (.I(\register_file[29][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13372__A2 (.I(\register_file[29][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__A2 (.I(\register_file[29][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13374__A2 (.I(\register_file[29][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A2 (.I(\register_file[29][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A2 (.I(\register_file[29][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__A2 (.I(\register_file[29][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A2 (.I(\register_file[29][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A2 (.I(\register_file[29][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13379__A2 (.I(\register_file[29][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A2 (.I(\register_file[29][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A2 (.I(\register_file[29][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13381__A2 (.I(\register_file[29][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A2 (.I(\register_file[29][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(\register_file[29][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13383__A2 (.I(\register_file[29][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A2 (.I(\register_file[29][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A2 (.I(\register_file[29][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__A2 (.I(\register_file[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13320__A2 (.I(\register_file[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A2 (.I(\register_file[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13387__A2 (.I(\register_file[29][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__A2 (.I(\register_file[29][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A2 (.I(\register_file[29][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__A2 (.I(\register_file[29][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A2 (.I(\register_file[29][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__I (.I(\register_file[29][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13894__A2 (.I(\register_file[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13323__A2 (.I(\register_file[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(\register_file[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13959__A2 (.I(\register_file[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13325__A2 (.I(\register_file[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A2 (.I(\register_file[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14049__A2 (.I(\register_file[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13329__A2 (.I(\register_file[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A2 (.I(\register_file[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14131__A2 (.I(\register_file[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13331__A2 (.I(\register_file[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A2 (.I(\register_file[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14307__A2 (.I(\register_file[29][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A2 (.I(\register_file[29][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(\register_file[29][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14390__A2 (.I(\register_file[29][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13338__A2 (.I(\register_file[29][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A2 (.I(\register_file[29][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14535__A2 (.I(\register_file[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A2 (.I(\register_file[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A2 (.I(\register_file[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14622__A2 (.I(\register_file[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A2 (.I(\register_file[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A2 (.I(\register_file[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14704__A2 (.I(\register_file[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(\register_file[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A2 (.I(\register_file[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14790__A2 (.I(\register_file[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A2 (.I(\register_file[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A2 (.I(\register_file[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14873__A2 (.I(\register_file[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A2 (.I(\register_file[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A2 (.I(\register_file[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14957__A2 (.I(\register_file[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A2 (.I(\register_file[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A2 (.I(\register_file[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15044__A2 (.I(\register_file[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A2 (.I(\register_file[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A2 (.I(\register_file[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15126__A2 (.I(\register_file[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A2 (.I(\register_file[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A2 (.I(\register_file[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15210__A2 (.I(\register_file[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A2 (.I(\register_file[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A2 (.I(\register_file[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15293__A2 (.I(\register_file[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A2 (.I(\register_file[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A2 (.I(\register_file[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15377__A2 (.I(\register_file[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A2 (.I(\register_file[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A2 (.I(\register_file[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15465__A2 (.I(\register_file[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A2 (.I(\register_file[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A2 (.I(\register_file[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15548__A2 (.I(\register_file[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A2 (.I(\register_file[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A2 (.I(\register_file[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A2 (.I(\register_file[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A2 (.I(\register_file[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A2 (.I(\register_file[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A2 (.I(\register_file[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A2 (.I(\register_file[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(\register_file[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A2 (.I(\register_file[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A2 (.I(\register_file[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A2 (.I(\register_file[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A2 (.I(\register_file[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A2 (.I(\register_file[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A2 (.I(\register_file[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A2 (.I(\register_file[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A2 (.I(\register_file[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A2 (.I(\register_file[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A2 (.I(\register_file[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A2 (.I(\register_file[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A2 (.I(\register_file[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13935__A2 (.I(\register_file[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__A2 (.I(\register_file[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A2 (.I(\register_file[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14023__A2 (.I(\register_file[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A2 (.I(\register_file[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A2 (.I(\register_file[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14108__A2 (.I(\register_file[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A2 (.I(\register_file[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A2 (.I(\register_file[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14282__A2 (.I(\register_file[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A2 (.I(\register_file[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(\register_file[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14368__A2 (.I(\register_file[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A2 (.I(\register_file[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(\register_file[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14451__A2 (.I(\register_file[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A2 (.I(\register_file[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A2 (.I(\register_file[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14478__A2 (.I(\register_file[30][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A2 (.I(\register_file[30][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A2 (.I(\register_file[30][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14560__A2 (.I(\register_file[30][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A2 (.I(\register_file[30][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A2 (.I(\register_file[30][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14644__A2 (.I(\register_file[30][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A2 (.I(\register_file[30][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A2 (.I(\register_file[30][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14731__A2 (.I(\register_file[30][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A2 (.I(\register_file[30][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A2 (.I(\register_file[30][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14815__A2 (.I(\register_file[30][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__A2 (.I(\register_file[30][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A2 (.I(\register_file[30][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14982__A2 (.I(\register_file[30][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(\register_file[30][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A2 (.I(\register_file[30][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15066__A2 (.I(\register_file[30][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A2 (.I(\register_file[30][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A2 (.I(\register_file[30][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15320__A2 (.I(\register_file[30][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A2 (.I(\register_file[30][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A2 (.I(\register_file[30][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15421__A2 (.I(\register_file[30][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A2 (.I(\register_file[30][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A2 (.I(\register_file[30][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15509__A2 (.I(\register_file[30][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A2 (.I(\register_file[30][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A2 (.I(\register_file[30][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15574__A2 (.I(\register_file[30][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__A2 (.I(\register_file[30][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A2 (.I(\register_file[30][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A2 (.I(\register_file[30][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A2 (.I(\register_file[30][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A2 (.I(\register_file[30][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__A2 (.I(\register_file[30][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A2 (.I(\register_file[30][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A2 (.I(\register_file[30][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A2 (.I(\register_file[30][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A2 (.I(\register_file[30][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A2 (.I(\register_file[30][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A2 (.I(\register_file[30][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__A2 (.I(\register_file[30][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A2 (.I(\register_file[30][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A2 (.I(\register_file[30][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A2 (.I(\register_file[30][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A2 (.I(\register_file[30][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13896__A2 (.I(\register_file[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A2 (.I(\register_file[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(\register_file[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13962__A2 (.I(\register_file[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A2 (.I(\register_file[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A2 (.I(\register_file[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14051__A2 (.I(\register_file[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A2 (.I(\register_file[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A2 (.I(\register_file[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14133__A2 (.I(\register_file[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A2 (.I(\register_file[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(\register_file[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14221__A2 (.I(\register_file[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A2 (.I(\register_file[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(\register_file[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14309__A2 (.I(\register_file[30][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A2 (.I(\register_file[30][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(\register_file[30][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14393__A2 (.I(\register_file[30][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__A2 (.I(\register_file[30][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A2 (.I(\register_file[30][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14479__A2 (.I(\register_file[31][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12216__A2 (.I(\register_file[31][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A2 (.I(\register_file[31][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14562__A2 (.I(\register_file[31][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12219__A2 (.I(\register_file[31][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A2 (.I(\register_file[31][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14645__A2 (.I(\register_file[31][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12222__A2 (.I(\register_file[31][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A2 (.I(\register_file[31][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14732__A2 (.I(\register_file[31][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12226__A2 (.I(\register_file[31][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A2 (.I(\register_file[31][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14817__A2 (.I(\register_file[31][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__A2 (.I(\register_file[31][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A2 (.I(\register_file[31][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14901__A2 (.I(\register_file[31][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__A2 (.I(\register_file[31][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(\register_file[31][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14984__A2 (.I(\register_file[31][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12236__A2 (.I(\register_file[31][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A2 (.I(\register_file[31][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15067__A2 (.I(\register_file[31][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__A2 (.I(\register_file[31][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A2 (.I(\register_file[31][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15174__A2 (.I(\register_file[31][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12243__A2 (.I(\register_file[31][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A2 (.I(\register_file[31][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15256__A2 (.I(\register_file[31][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12246__A2 (.I(\register_file[31][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A2 (.I(\register_file[31][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15321__A2 (.I(\register_file[31][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12250__A2 (.I(\register_file[31][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__A2 (.I(\register_file[31][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15422__A2 (.I(\register_file[31][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12253__A2 (.I(\register_file[31][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A2 (.I(\register_file[31][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15512__A2 (.I(\register_file[31][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12256__A2 (.I(\register_file[31][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(\register_file[31][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15575__A2 (.I(\register_file[31][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12260__A2 (.I(\register_file[31][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A2 (.I(\register_file[31][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12263__A2 (.I(\register_file[31][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A2 (.I(\register_file[31][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A2 (.I(\register_file[31][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12267__A2 (.I(\register_file[31][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A2 (.I(\register_file[31][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A2 (.I(\register_file[31][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12270__A2 (.I(\register_file[31][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A2 (.I(\register_file[31][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(\register_file[31][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12273__A2 (.I(\register_file[31][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__A2 (.I(\register_file[31][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A2 (.I(\register_file[31][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12276__A2 (.I(\register_file[31][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__A2 (.I(\register_file[31][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A2 (.I(\register_file[31][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12279__A2 (.I(\register_file[31][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A2 (.I(\register_file[31][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A2 (.I(\register_file[31][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12282__A2 (.I(\register_file[31][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A2 (.I(\register_file[31][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A2 (.I(\register_file[31][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12285__A2 (.I(\register_file[31][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A2 (.I(\register_file[31][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__I (.I(\register_file[31][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13897__A2 (.I(\register_file[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12191__A2 (.I(\register_file[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A2 (.I(\register_file[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14052__A2 (.I(\register_file[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12199__A2 (.I(\register_file[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A2 (.I(\register_file[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14136__A2 (.I(\register_file[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12202__A2 (.I(\register_file[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A2 (.I(\register_file[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14222__A2 (.I(\register_file[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12205__A2 (.I(\register_file[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A2 (.I(\register_file[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14310__A2 (.I(\register_file[31][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A2 (.I(\register_file[31][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A2 (.I(\register_file[31][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14395__A2 (.I(\register_file[31][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12212__A2 (.I(\register_file[31][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A2 (.I(\register_file[31][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13660__I (.I(\register_file[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12100__A2 (.I(\register_file[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A2 (.I(\register_file[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14623__I (.I(\register_file[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12127__A2 (.I(\register_file[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A2 (.I(\register_file[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14705__I (.I(\register_file[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12129__A2 (.I(\register_file[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A2 (.I(\register_file[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15127__I (.I(\register_file[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12141__A2 (.I(\register_file[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A2 (.I(\register_file[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15378__I (.I(\register_file[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__A2 (.I(\register_file[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A2 (.I(\register_file[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15466__I (.I(\register_file[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12151__A2 (.I(\register_file[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A2 (.I(\register_file[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15549__I (.I(\register_file[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__A2 (.I(\register_file[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A2 (.I(\register_file[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12156__A2 (.I(\register_file[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A2 (.I(\register_file[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__I (.I(\register_file[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12167__A2 (.I(\register_file[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A2 (.I(\register_file[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__I (.I(\register_file[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12169__A2 (.I(\register_file[3][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A2 (.I(\register_file[3][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__I (.I(\register_file[3][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13847__I (.I(\register_file[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__A2 (.I(\register_file[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A2 (.I(\register_file[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12171__A2 (.I(\register_file[3][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A2 (.I(\register_file[3][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__I (.I(\register_file[3][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12173__A2 (.I(\register_file[3][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A2 (.I(\register_file[3][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A2 (.I(\register_file[3][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13936__I (.I(\register_file[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__A2 (.I(\register_file[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A2 (.I(\register_file[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14024__I (.I(\register_file[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12109__A2 (.I(\register_file[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A2 (.I(\register_file[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14109__I (.I(\register_file[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12113__A2 (.I(\register_file[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A2 (.I(\register_file[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14200__I (.I(\register_file[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12115__A2 (.I(\register_file[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A2 (.I(\register_file[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14283__I (.I(\register_file[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__A2 (.I(\register_file[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A2 (.I(\register_file[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14369__I (.I(\register_file[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12120__A2 (.I(\register_file[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A2 (.I(\register_file[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14612__I (.I(\register_file[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A2 (.I(\register_file[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15203__I (.I(\register_file[4][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A2 (.I(\register_file[4][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15285__I (.I(\register_file[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A2 (.I(\register_file[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13748__I (.I(\register_file[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A2 (.I(\register_file[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15455__I (.I(\register_file[4][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A2 (.I(\register_file[4][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A2 (.I(\register_file[4][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__I (.I(\register_file[4][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A2 (.I(\register_file[4][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__I (.I(\register_file[4][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__A2 (.I(\register_file[4][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__I (.I(\register_file[4][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A2 (.I(\register_file[4][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__I (.I(\register_file[4][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14100__I (.I(\register_file[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A2 (.I(\register_file[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14275__I (.I(\register_file[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(\register_file[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14614__I (.I(\register_file[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11967__A2 (.I(\register_file[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A2 (.I(\register_file[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14699__I (.I(\register_file[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__A2 (.I(\register_file[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A2 (.I(\register_file[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15205__I (.I(\register_file[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11984__A2 (.I(\register_file[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A2 (.I(\register_file[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15287__I (.I(\register_file[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11986__A2 (.I(\register_file[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A2 (.I(\register_file[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13750__I (.I(\register_file[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11942__A2 (.I(\register_file[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A2 (.I(\register_file[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15371__I (.I(\register_file[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__A2 (.I(\register_file[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A2 (.I(\register_file[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15457__I (.I(\register_file[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11991__A2 (.I(\register_file[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A2 (.I(\register_file[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15543__I (.I(\register_file[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__A2 (.I(\register_file[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A2 (.I(\register_file[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12003__A2 (.I(\register_file[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A2 (.I(\register_file[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__I (.I(\register_file[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__A2 (.I(\register_file[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A2 (.I(\register_file[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__I (.I(\register_file[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__A2 (.I(\register_file[5][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A2 (.I(\register_file[5][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__I (.I(\register_file[5][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13930__I (.I(\register_file[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11947__A2 (.I(\register_file[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A2 (.I(\register_file[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14102__I (.I(\register_file[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__A2 (.I(\register_file[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A2 (.I(\register_file[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14277__I (.I(\register_file[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__A2 (.I(\register_file[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A2 (.I(\register_file[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14363__I (.I(\register_file[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__A2 (.I(\register_file[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A2 (.I(\register_file[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14445__I (.I(\register_file[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__A2 (.I(\register_file[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A2 (.I(\register_file[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14607__A2 (.I(\register_file[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11887__A2 (.I(\register_file[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(\register_file[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15199__A2 (.I(\register_file[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11904__A2 (.I(\register_file[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A2 (.I(\register_file[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15365__A2 (.I(\register_file[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__A2 (.I(\register_file[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A2 (.I(\register_file[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15450__A2 (.I(\register_file[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11911__A2 (.I(\register_file[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A2 (.I(\register_file[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15536__A2 (.I(\register_file[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__A2 (.I(\register_file[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A2 (.I(\register_file[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11916__A2 (.I(\register_file[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A2 (.I(\register_file[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A2 (.I(\register_file[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11918__A2 (.I(\register_file[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A2 (.I(\register_file[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A2 (.I(\register_file[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11923__A2 (.I(\register_file[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A2 (.I(\register_file[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A2 (.I(\register_file[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11927__A2 (.I(\register_file[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A2 (.I(\register_file[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A2 (.I(\register_file[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__A2 (.I(\register_file[6][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__A2 (.I(\register_file[6][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A2 (.I(\register_file[6][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13924__A2 (.I(\register_file[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11867__A2 (.I(\register_file[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A2 (.I(\register_file[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14009__A2 (.I(\register_file[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11869__A2 (.I(\register_file[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A2 (.I(\register_file[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14096__A2 (.I(\register_file[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11873__A2 (.I(\register_file[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A2 (.I(\register_file[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14184__A2 (.I(\register_file[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11875__A2 (.I(\register_file[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A2 (.I(\register_file[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14270__A2 (.I(\register_file[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__A2 (.I(\register_file[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A2 (.I(\register_file[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14357__A2 (.I(\register_file[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11880__A2 (.I(\register_file[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A2 (.I(\register_file[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14608__I (.I(\register_file[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__A2 (.I(\register_file[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A2 (.I(\register_file[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14693__I (.I(\register_file[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11809__A2 (.I(\register_file[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A2 (.I(\register_file[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14861__I (.I(\register_file[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__A2 (.I(\register_file[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A2 (.I(\register_file[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15030__I (.I(\register_file[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__A2 (.I(\register_file[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A2 (.I(\register_file[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15115__I (.I(\register_file[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11821__A2 (.I(\register_file[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A2 (.I(\register_file[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15200__I (.I(\register_file[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11824__A2 (.I(\register_file[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A2 (.I(\register_file[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13744__I (.I(\register_file[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__A2 (.I(\register_file[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A2 (.I(\register_file[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15366__I (.I(\register_file[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11829__A2 (.I(\register_file[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A2 (.I(\register_file[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15451__I (.I(\register_file[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__A2 (.I(\register_file[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A2 (.I(\register_file[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15537__I (.I(\register_file[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__A2 (.I(\register_file[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A2 (.I(\register_file[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__A2 (.I(\register_file[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A2 (.I(\register_file[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__I (.I(\register_file[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11843__A2 (.I(\register_file[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A2 (.I(\register_file[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__I (.I(\register_file[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11847__A2 (.I(\register_file[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A2 (.I(\register_file[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__I (.I(\register_file[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11849__A2 (.I(\register_file[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A2 (.I(\register_file[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__I (.I(\register_file[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14010__I (.I(\register_file[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11789__A2 (.I(\register_file[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A2 (.I(\register_file[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14097__I (.I(\register_file[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__A2 (.I(\register_file[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A2 (.I(\register_file[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14185__I (.I(\register_file[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11795__A2 (.I(\register_file[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(\register_file[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14271__I (.I(\register_file[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11797__A2 (.I(\register_file[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A2 (.I(\register_file[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14358__I (.I(\register_file[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__A2 (.I(\register_file[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A2 (.I(\register_file[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14439__I (.I(\register_file[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11802__A2 (.I(\register_file[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A2 (.I(\register_file[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__A2 (.I(\register_file[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__A2 (.I(\register_file[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A2 (.I(\register_file[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14585__A2 (.I(\register_file[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__A2 (.I(\register_file[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A2 (.I(\register_file[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14673__A2 (.I(\register_file[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11710__A2 (.I(\register_file[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A2 (.I(\register_file[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14759__A2 (.I(\register_file[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A2 (.I(\register_file[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A2 (.I(\register_file[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14843__A2 (.I(\register_file[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__A2 (.I(\register_file[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A2 (.I(\register_file[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14924__A2 (.I(\register_file[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__A2 (.I(\register_file[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A2 (.I(\register_file[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15007__A2 (.I(\register_file[8][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11724__A2 (.I(\register_file[8][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A2 (.I(\register_file[8][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15095__A2 (.I(\register_file[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__A2 (.I(\register_file[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A2 (.I(\register_file[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15179__A2 (.I(\register_file[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__A2 (.I(\register_file[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A2 (.I(\register_file[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13721__A2 (.I(\register_file[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__A2 (.I(\register_file[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A2 (.I(\register_file[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15344__A2 (.I(\register_file[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11738__A2 (.I(\register_file[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A2 (.I(\register_file[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15428__A2 (.I(\register_file[8][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__A2 (.I(\register_file[8][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A2 (.I(\register_file[8][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15517__A2 (.I(\register_file[8][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11744__A2 (.I(\register_file[8][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A2 (.I(\register_file[8][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15601__A2 (.I(\register_file[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__A2 (.I(\register_file[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(\register_file[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11751__A2 (.I(\register_file[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__A2 (.I(\register_file[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A2 (.I(\register_file[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11755__A2 (.I(\register_file[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A2 (.I(\register_file[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A2 (.I(\register_file[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__A2 (.I(\register_file[8][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A2 (.I(\register_file[8][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(\register_file[8][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__A2 (.I(\register_file[8][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A2 (.I(\register_file[8][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A2 (.I(\register_file[8][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__A2 (.I(\register_file[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A2 (.I(\register_file[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A2 (.I(\register_file[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11767__A2 (.I(\register_file[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A2 (.I(\register_file[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A2 (.I(\register_file[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13814__A2 (.I(\register_file[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__A2 (.I(\register_file[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A2 (.I(\register_file[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__A2 (.I(\register_file[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A2 (.I(\register_file[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A2 (.I(\register_file[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__A2 (.I(\register_file[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A2 (.I(\register_file[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A2 (.I(\register_file[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13902__A2 (.I(\register_file[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__A2 (.I(\register_file[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A2 (.I(\register_file[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13992__A2 (.I(\register_file[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__A2 (.I(\register_file[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A2 (.I(\register_file[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14075__A2 (.I(\register_file[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__A2 (.I(\register_file[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A2 (.I(\register_file[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14160__A2 (.I(\register_file[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11690__A2 (.I(\register_file[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(\register_file[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14250__A2 (.I(\register_file[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__A2 (.I(\register_file[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A2 (.I(\register_file[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14337__A2 (.I(\register_file[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__A2 (.I(\register_file[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(\register_file[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14421__A2 (.I(\register_file[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__A2 (.I(\register_file[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A2 (.I(\register_file[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14587__A2 (.I(\register_file[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13423__A2 (.I(\register_file[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A2 (.I(\register_file[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14925__A2 (.I(\register_file[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13433__A2 (.I(\register_file[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(\register_file[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13723__A2 (.I(\register_file[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13398__A2 (.I(\register_file[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A2 (.I(\register_file[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15345__A2 (.I(\register_file[9][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13445__A2 (.I(\register_file[9][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A2 (.I(\register_file[9][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15430__A2 (.I(\register_file[9][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13447__A2 (.I(\register_file[9][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A2 (.I(\register_file[9][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15518__A2 (.I(\register_file[9][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13449__A2 (.I(\register_file[9][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A2 (.I(\register_file[9][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15602__A2 (.I(\register_file[9][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13452__A2 (.I(\register_file[9][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A2 (.I(\register_file[9][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13454__A2 (.I(\register_file[9][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A2 (.I(\register_file[9][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A2 (.I(\register_file[9][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13457__A2 (.I(\register_file[9][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A2 (.I(\register_file[9][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A2 (.I(\register_file[9][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13459__A2 (.I(\register_file[9][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A2 (.I(\register_file[9][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A2 (.I(\register_file[9][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13461__A2 (.I(\register_file[9][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A2 (.I(\register_file[9][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A2 (.I(\register_file[9][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13465__A2 (.I(\register_file[9][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A2 (.I(\register_file[9][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A2 (.I(\register_file[9][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13815__A2 (.I(\register_file[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13400__A2 (.I(\register_file[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A2 (.I(\register_file[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13467__A2 (.I(\register_file[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A2 (.I(\register_file[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(\register_file[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13903__A2 (.I(\register_file[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13403__A2 (.I(\register_file[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A2 (.I(\register_file[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13993__A2 (.I(\register_file[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13405__A2 (.I(\register_file[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(\register_file[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14076__A2 (.I(\register_file[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13409__A2 (.I(\register_file[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A2 (.I(\register_file[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14162__A2 (.I(\register_file[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13411__A2 (.I(\register_file[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A2 (.I(\register_file[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14338__A2 (.I(\register_file[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13416__A2 (.I(\register_file[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(\register_file[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14422__A2 (.I(\register_file[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13418__A2 (.I(\register_file[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A2 (.I(\register_file[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A3 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A3 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A3 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13476__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13471__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13502__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13482__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13500__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13482__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13908__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13666__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13544__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13487__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13988__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13672__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13583__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12049__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12052__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12054__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12057__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12059__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12061__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12064__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12066__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12022__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__A2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12083__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12087__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12089__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12024__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12091__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12093__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__A2 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12033__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12042__A2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output74_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output80_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output81_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output82_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output83_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output84_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output85_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output86_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output87_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output88_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output89_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output90_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output91_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16031__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15999__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16000__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16001__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16002__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16003__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16512__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15967__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16032__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15936__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16447__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16448__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16511__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16352__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16351__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15648__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15647__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16096__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15935__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16095__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16543__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15938__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15937__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15743__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15744__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16576__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16575__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15840__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16544__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15871__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15903__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15808__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16191__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15807__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16192__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15776__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16579__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15839__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16098__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16099__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16097__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15939__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16577__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16578__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15711__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16319__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16416__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15712__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16383__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16415__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16159__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16384__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16287__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16545__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16547__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16127__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16128__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16546__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15682__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15681__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15617__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15679__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15615__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15616__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16320__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15649__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15619__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15683__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15618__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16514__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16515__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15841__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16481__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16513__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15873__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16224__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15905__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15678__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15614__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16255__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16223__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16158__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16382__CLK (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16381__CLK (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15774__CLK (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16317__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16285__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16318__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16222__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16190__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16126__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16189__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16125__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16221__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16253__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16157__CLK (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16156__CLK (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16188__CLK (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15708__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15676__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16105__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15945__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16106__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15847__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15878__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16520__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16487__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16488__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16486__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16518__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16519__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15810__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15942__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16583__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16582__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15811__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15809__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15874__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15907__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15875__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16450__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15842__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16483__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15777__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15778__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15713__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15745__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15746__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15651__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16482__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16101__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16100__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15747__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15715__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16449__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15714__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15843__CLK (.I(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15779__CLK (.I(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16451__CLK (.I(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16354__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16355__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16353__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15940__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16385__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16419__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16417__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16418__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16516__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16517__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16130__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16322__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16387__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16386__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16485__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15844__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15845__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16131__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15908__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15812__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15876__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16162__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16549__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16161__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16163__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16321__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16129__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16452__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16453__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15717__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15749__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15653__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15652__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15748__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16548__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16194__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16193__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15716__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15684__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16257__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16258__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16195__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15620__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15621__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15685__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16226__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16225__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16421__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16324__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16420__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16389__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16292__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16356__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16357__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16261__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16164__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16260__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16293__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16388__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16229__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16227__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16259__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16133__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16328__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16327__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16294__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16296__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16295__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16165__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16197__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16230__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16360__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16358__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16359__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16390__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16392__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16391__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15750__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15686__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16424__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16422__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16552__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15687__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16551__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16550__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15623__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15719__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15654__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15655__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15720__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15718__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16200__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16168__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16167__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16199__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16135__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16232__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16138__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16169__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16170__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15658__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15721__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15657__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15656__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16361__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16265__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16266__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16362__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16201__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16202__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16203__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16298__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16297__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16394__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16393__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16234__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16426__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16139__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16171__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16204__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16425__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15626__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15627__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16330__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16329__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15753__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15690__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15625__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15814__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15815__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15816__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15879__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15880__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15912__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15911__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15910__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15913__CLK (.I(clknet_leaf_111_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15850__CLK (.I(clknet_leaf_111_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15849__CLK (.I(clknet_leaf_111_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15882__CLK (.I(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15914__CLK (.I(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15915__CLK (.I(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16585__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16490__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15947__CLK (.I(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16587__CLK (.I(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16586__CLK (.I(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16589__CLK (.I(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15949__CLK (.I(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15948__CLK (.I(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15916__CLK (.I(clknet_leaf_122_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15852__CLK (.I(clknet_leaf_122_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15851__CLK (.I(clknet_leaf_122_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16524__CLK (.I(clknet_leaf_123_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15789__CLK (.I(clknet_leaf_123_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15788__CLK (.I(clknet_leaf_123_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16526__CLK (.I(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16525__CLK (.I(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16493__CLK (.I(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15854__CLK (.I(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15853__CLK (.I(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16527__CLK (.I(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15790__CLK (.I(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15823__CLK (.I(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15791__CLK (.I(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15855__CLK (.I(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15628__CLK (.I(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15629__CLK (.I(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15691__CLK (.I(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15660__CLK (.I(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16235__CLK (.I(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15755__CLK (.I(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15756__CLK (.I(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15723__CLK (.I(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15725__CLK (.I(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16205__CLK (.I(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16299__CLK (.I(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16173__CLK (.I(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16268__CLK (.I(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16267__CLK (.I(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16172__CLK (.I(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16395__CLK (.I(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16300__CLK (.I(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16269__CLK (.I(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16140__CLK (.I(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16237__CLK (.I(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16141__CLK (.I(clknet_leaf_140_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16428__CLK (.I(clknet_leaf_140_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16363__CLK (.I(clknet_leaf_140_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16396__CLK (.I(clknet_leaf_140_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16364__CLK (.I(clknet_leaf_140_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16397__CLK (.I(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16429__CLK (.I(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16333__CLK (.I(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15661__CLK (.I(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16398__CLK (.I(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16367__CLK (.I(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16175__CLK (.I(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16366__CLK (.I(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16399__CLK (.I(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16431__CLK (.I(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16334__CLK (.I(clknet_leaf_145_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16238__CLK (.I(clknet_leaf_145_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16303__CLK (.I(clknet_leaf_145_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16302__CLK (.I(clknet_leaf_145_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15663__CLK (.I(clknet_leaf_146_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15759__CLK (.I(clknet_leaf_146_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15726__CLK (.I(clknet_leaf_146_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16335__CLK (.I(clknet_leaf_146_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16463__CLK (.I(clknet_leaf_148_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15758__CLK (.I(clknet_leaf_148_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15693__CLK (.I(clknet_leaf_148_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15757__CLK (.I(clknet_leaf_148_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16559__CLK (.I(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16558__CLK (.I(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15822__CLK (.I(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16240__CLK (.I(clknet_leaf_151_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16148__CLK (.I(clknet_leaf_151_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16147__CLK (.I(clknet_leaf_151_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15631__CLK (.I(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15695__CLK (.I(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15694__CLK (.I(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15630__CLK (.I(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16270__CLK (.I(clknet_leaf_153_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16143__CLK (.I(clknet_leaf_153_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16142__CLK (.I(clknet_leaf_153_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16239__CLK (.I(clknet_leaf_153_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16241__CLK (.I(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16242__CLK (.I(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16144__CLK (.I(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16145__CLK (.I(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16146__CLK (.I(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16337__CLK (.I(clknet_leaf_157_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16211__CLK (.I(clknet_leaf_157_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16212__CLK (.I(clknet_leaf_157_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16273__CLK (.I(clknet_leaf_158_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16306__CLK (.I(clknet_leaf_158_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16274__CLK (.I(clknet_leaf_158_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16304__CLK (.I(clknet_leaf_158_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16370__CLK (.I(clknet_leaf_159_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16305__CLK (.I(clknet_leaf_159_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16402__CLK (.I(clknet_leaf_159_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16400__CLK (.I(clknet_leaf_160_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16401__CLK (.I(clknet_leaf_160_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16369__CLK (.I(clknet_leaf_160_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16336__CLK (.I(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16180__CLK (.I(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16338__CLK (.I(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16433__CLK (.I(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16561__CLK (.I(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15633__CLK (.I(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15696__CLK (.I(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15632__CLK (.I(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16434__CLK (.I(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15729__CLK (.I(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16464__CLK (.I(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16466__CLK (.I(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15728__CLK (.I(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15697__CLK (.I(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16436__CLK (.I(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16435__CLK (.I(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16467__CLK (.I(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16468__CLK (.I(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15824__CLK (.I(clknet_leaf_169_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15792__CLK (.I(clknet_leaf_169_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15826__CLK (.I(clknet_leaf_169_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15858__CLK (.I(clknet_leaf_171_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15890__CLK (.I(clknet_leaf_171_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15889__CLK (.I(clknet_leaf_171_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15857__CLK (.I(clknet_leaf_171_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16529__CLK (.I(clknet_leaf_172_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15795__CLK (.I(clknet_leaf_172_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15796__CLK (.I(clknet_leaf_172_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15828__CLK (.I(clknet_leaf_172_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16528__CLK (.I(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15664__CLK (.I(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15665__CLK (.I(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15761__CLK (.I(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15760__CLK (.I(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15730__CLK (.I(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16404__CLK (.I(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15827__CLK (.I(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16500__CLK (.I(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16499__CLK (.I(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16496__CLK (.I(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16532__CLK (.I(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16531__CLK (.I(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15860__CLK (.I(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16530__CLK (.I(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16498__CLK (.I(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16497__CLK (.I(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16592__CLK (.I(clknet_leaf_176_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15859__CLK (.I(clknet_leaf_176_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16594__CLK (.I(clknet_leaf_176_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15732__CLK (.I(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15731__CLK (.I(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15763__CLK (.I(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15764__CLK (.I(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15762__CLK (.I(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15635__CLK (.I(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15634__CLK (.I(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15698__CLK (.I(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15666__CLK (.I(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16593__CLK (.I(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16150__CLK (.I(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16149__CLK (.I(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16243__CLK (.I(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16244__CLK (.I(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15919__CLK (.I(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15888__CLK (.I(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15920__CLK (.I(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15887__CLK (.I(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15886__CLK (.I(clknet_leaf_187_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15918__CLK (.I(clknet_leaf_187_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16494__CLK (.I(clknet_leaf_188_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16495__CLK (.I(clknet_leaf_188_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16590__CLK (.I(clknet_leaf_188_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15950__CLK (.I(clknet_leaf_189_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15951__CLK (.I(clknet_leaf_189_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16591__CLK (.I(clknet_leaf_189_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16152__CLK (.I(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16151__CLK (.I(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16183__CLK (.I(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16247__CLK (.I(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16111__CLK (.I(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16153__CLK (.I(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16280__CLK (.I(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16184__CLK (.I(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16249__CLK (.I(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16281__CLK (.I(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16248__CLK (.I(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16108__CLK (.I(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16107__CLK (.I(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16344__CLK (.I(clknet_leaf_195_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16408__CLK (.I(clknet_leaf_195_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16216__CLK (.I(clknet_leaf_196_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16185__CLK (.I(clknet_leaf_196_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16217__CLK (.I(clknet_leaf_196_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16345__CLK (.I(clknet_leaf_196_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15704__CLK (.I(clknet_leaf_196_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16343__CLK (.I(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16215__CLK (.I(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16279__CLK (.I(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15640__CLK (.I(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15736__CLK (.I(clknet_leaf_199_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15705__CLK (.I(clknet_leaf_199_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15641__CLK (.I(clknet_leaf_199_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16377__CLK (.I(clknet_leaf_202_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16375__CLK (.I(clknet_leaf_202_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16473__CLK (.I(clknet_leaf_202_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16438__CLK (.I(clknet_leaf_204_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16439__CLK (.I(clknet_leaf_204_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16440__CLK (.I(clknet_leaf_204_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15798__CLK (.I(clknet_leaf_204_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15797__CLK (.I(clknet_leaf_205_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16437__CLK (.I(clknet_leaf_205_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16214__CLK (.I(clknet_leaf_207_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16278__CLK (.I(clknet_leaf_207_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16372__CLK (.I(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16275__CLK (.I(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16307__CLK (.I(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15924__CLK (.I(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15667__CLK (.I(clknet_leaf_210_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15668__CLK (.I(clknet_leaf_210_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15636__CLK (.I(clknet_leaf_210_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16339__CLK (.I(clknet_leaf_210_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16564__CLK (.I(clknet_leaf_210_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16371__CLK (.I(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15733__CLK (.I(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15701__CLK (.I(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15637__CLK (.I(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16405__CLK (.I(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15923__CLK (.I(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15891__CLK (.I(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15892__CLK (.I(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16595__CLK (.I(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16406__CLK (.I(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16596__CLK (.I(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15799__CLK (.I(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16469__CLK (.I(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16471__CLK (.I(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16567__CLK (.I(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16565__CLK (.I(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16566__CLK (.I(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15953__CLK (.I(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15954__CLK (.I(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15952__CLK (.I(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15893__CLK (.I(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16470__CLK (.I(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16116__CLK (.I(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15956__CLK (.I(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15957__CLK (.I(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16117__CLK (.I(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15671__CLK (.I(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15669__CLK (.I(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16598__CLK (.I(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15767__CLK (.I(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15766__CLK (.I(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15955__CLK (.I(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16112__CLK (.I(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16113__CLK (.I(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16535__CLK (.I(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16534__CLK (.I(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15985__CLK (.I(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15986__CLK (.I(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15988__CLK (.I(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16016__CLK (.I(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16018__CLK (.I(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16017__CLK (.I(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16114__CLK (.I(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16084__CLK (.I(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16050__CLK (.I(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16048__CLK (.I(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16049__CLK (.I(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16052__CLK (.I(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15984__CLK (.I(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16082__CLK (.I(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16051__CLK (.I(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16083__CLK (.I(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16085__CLK (.I(clknet_leaf_233_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16053__CLK (.I(clknet_leaf_233_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15989__CLK (.I(clknet_leaf_233_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16079__CLK (.I(clknet_leaf_234_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16087__CLK (.I(clknet_leaf_234_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16054__CLK (.I(clknet_leaf_234_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16086__CLK (.I(clknet_leaf_234_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16080__CLK (.I(clknet_leaf_234_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16118__CLK (.I(clknet_leaf_238_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16021__CLK (.I(clknet_leaf_238_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15672__CLK (.I(clknet_leaf_240_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16376__CLK (.I(clknet_leaf_240_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16536__CLK (.I(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16537__CLK (.I(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16120__CLK (.I(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16121__CLK (.I(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15673__CLK (.I(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16024__CLK (.I(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16025__CLK (.I(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15993__CLK (.I(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16015__CLK (.I(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15992__CLK (.I(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16056__CLK (.I(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15983__CLK (.I(clknet_leaf_245_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15982__CLK (.I(clknet_leaf_245_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16046__CLK (.I(clknet_leaf_245_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16047__CLK (.I(clknet_leaf_245_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16058__CLK (.I(clknet_leaf_248_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16090__CLK (.I(clknet_leaf_248_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16089__CLK (.I(clknet_leaf_248_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16026__CLK (.I(clknet_leaf_252_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15994__CLK (.I(clknet_leaf_252_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16027__CLK (.I(clknet_leaf_252_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16122__CLK (.I(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16570__CLK (.I(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16602__CLK (.I(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16474__CLK (.I(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15962__CLK (.I(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15770__CLK (.I(clknet_leaf_255_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15866__CLK (.I(clknet_leaf_255_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16378__CLK (.I(clknet_leaf_255_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15961__CLK (.I(clknet_leaf_257_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16601__CLK (.I(clknet_leaf_257_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16600__CLK (.I(clknet_leaf_257_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15674__CLK (.I(clknet_leaf_257_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15865__CLK (.I(clknet_leaf_260_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15832__CLK (.I(clknet_leaf_260_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15864__CLK (.I(clknet_leaf_260_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15801__CLK (.I(clknet_leaf_261_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15800__CLK (.I(clknet_leaf_261_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15897__CLK (.I(clknet_leaf_261_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15833__CLK (.I(clknet_leaf_263_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16569__CLK (.I(clknet_leaf_263_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16409__CLK (.I(clknet_leaf_263_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15834__CLK (.I(clknet_leaf_265_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15899__CLK (.I(clknet_leaf_265_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15931__CLK (.I(clknet_leaf_265_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15898__CLK (.I(clknet_leaf_265_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16251__CLK (.I(clknet_leaf_269_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16282__CLK (.I(clknet_leaf_269_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16250__CLK (.I(clknet_leaf_269_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16154__CLK (.I(clknet_leaf_269_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15643__CLK (.I(clknet_leaf_271_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15707__CLK (.I(clknet_leaf_271_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16380__CLK (.I(clknet_leaf_278_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16316__CLK (.I(clknet_leaf_278_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15805__CLK (.I(clknet_leaf_279_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15837__CLK (.I(clknet_leaf_279_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15836__CLK (.I(clknet_leaf_279_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15772__CLK (.I(clknet_leaf_279_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15644__CLK (.I(clknet_leaf_282_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16540__CLK (.I(clknet_leaf_282_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16476__CLK (.I(clknet_leaf_282_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15771__CLK (.I(clknet_leaf_283_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15900__CLK (.I(clknet_leaf_283_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15740__CLK (.I(clknet_leaf_283_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16603__CLK (.I(clknet_leaf_284_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15675__CLK (.I(clknet_leaf_284_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16379__CLK (.I(clknet_leaf_284_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16091__CLK (.I(clknet_leaf_288_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16059__CLK (.I(clknet_leaf_288_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15995__CLK (.I(clknet_leaf_288_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16123__CLK (.I(clknet_leaf_288_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16042__CLK (.I(clknet_leaf_289_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16073__CLK (.I(clknet_leaf_289_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16043__CLK (.I(clknet_leaf_289_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15978__CLK (.I(clknet_leaf_291_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15977__CLK (.I(clknet_leaf_291_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16041__CLK (.I(clknet_leaf_291_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15964__CLK (.I(clknet_leaf_293_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16028__CLK (.I(clknet_leaf_293_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16060__CLK (.I(clknet_leaf_293_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16039__CLK (.I(clknet_leaf_296_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16040__CLK (.I(clknet_leaf_296_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16008__CLK (.I(clknet_leaf_296_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16007__CLK (.I(clknet_leaf_297_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15976__CLK (.I(clknet_leaf_297_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15975__CLK (.I(clknet_leaf_297_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16509__CLK (.I(clknet_leaf_300_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16061__CLK (.I(clknet_leaf_300_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16062__CLK (.I(clknet_leaf_300_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16541__CLK (.I(clknet_leaf_301_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16477__CLK (.I(clknet_leaf_301_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16092__CLK (.I(clknet_leaf_301_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16349__CLK (.I(clknet_leaf_302_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15645__CLK (.I(clknet_leaf_302_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16542__CLK (.I(clknet_leaf_302_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16350__CLK (.I(clknet_leaf_303_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15902__CLK (.I(clknet_leaf_303_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16445__CLK (.I(clknet_leaf_304_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16446__CLK (.I(clknet_leaf_304_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15646__CLK (.I(clknet_leaf_304_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16573__CLK (.I(clknet_leaf_304_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16478__CLK (.I(clknet_leaf_305_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16510__CLK (.I(clknet_leaf_305_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16574__CLK (.I(clknet_leaf_305_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15934__CLK (.I(clknet_leaf_305_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15965__CLK (.I(clknet_leaf_307_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15997__CLK (.I(clknet_leaf_307_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15933__CLK (.I(clknet_leaf_307_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16070__CLK (.I(clknet_leaf_309_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16038__CLK (.I(clknet_leaf_309_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15974__CLK (.I(clknet_leaf_309_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16006__CLK (.I(clknet_leaf_309_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16069__CLK (.I(clknet_leaf_310_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16067__CLK (.I(clknet_leaf_310_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16066__CLK (.I(clknet_leaf_310_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15972__CLK (.I(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16005__CLK (.I(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15973__CLK (.I(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16065__CLK (.I(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16068__CLK (.I(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15970__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16004__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15971__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15969__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16035__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16033__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16034__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16037__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16036__CLK (.I(clknet_leaf_314_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_3__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_2__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_1__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_0__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_7__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_6__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_5__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_4__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_11__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_10__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_9__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_8__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_15__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_14__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_13__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_12__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_19__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_18__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_17__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_16__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_23__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_22__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_21__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_20__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_27__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_26__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_25__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_24__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_31__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_30__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_29__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_28__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_314_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_313_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15968__CLK (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16064__CLK (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_310_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_309_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15966__CLK (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_307_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_306_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_305_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_304_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_303_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16256__CLK (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15710__CLK (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15870__CLK (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_302_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_301_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_300_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_299_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_298_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_297_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_296_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_295_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15996__CLK (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_282_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_281_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_293_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_292_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_291_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16074__CLK (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_289_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_288_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_287_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_286_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_285_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_284_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_283_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_280_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_279_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_278_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16284__CLK (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_277_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_276_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_275_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_274_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15739__CLK (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_272_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_271_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_270_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_269_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15941__CLK (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15650__CLK (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15906__CLK (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16584__CLK (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15946__CLK (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15881__CLK (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15782__CLK (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16553__CLK (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16458__CLK (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_257_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_256_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_255_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_254_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_253_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_252_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_251_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_250_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_249_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_248_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16505__CLK (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_247_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_246_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_245_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_244_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_243_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_242_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_241_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_240_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15642__CLK (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_267_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16442__CLK (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_265_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_264_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_263_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_196_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_195_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_194_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_262_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_261_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_260_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_259_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_202_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_201_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16472__CLK (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_199_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16311__CLK (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_197_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_239_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_238_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_237_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16023__CLK (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_235_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_234_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_233_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_221_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_220_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16081__CLK (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_231_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_230_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_229_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_228_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16115__CLK (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_226_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_225_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_224_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_223_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_222_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_217_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_219_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_208_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_207_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_206_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_205_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_204_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_203_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_182_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_218_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_216_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_215_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_214_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_213_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_212_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_211_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_210_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_209_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_179_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_193_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16491__CLK (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16492__CLK (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16588__CLK (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_192_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_191_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_190_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_189_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_188_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_187_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_140_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_137_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_136_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15724__CLK (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15727__CLK (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_148_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_147_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_146_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_142_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16461__CLK (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_186_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_185_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16181__CLK (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_183_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_181_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_171_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_170_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_180_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_178_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_177_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_176_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_175_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_174_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_173_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_172_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_169_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_156_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_155_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_154_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_153_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_152_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_151_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_150_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_168_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_167_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_166_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_165_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_164_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16179__CLK (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_162_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_161_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_160_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_159_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_158_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_157_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1577 ();
endmodule

